`define BETA 00010011
`define BETA_WIDTH 8
`define BETA_INT_WIDTH 0
`define BETA_FRACT_WIDTH 8

`define DELTA_T 0000000011000101
`define DELTA_T_WIDTH 16
`define DELTA_T_INT_WIDTH 
`define DELTA_T_FRACT_WIDTH 16

`define ACC_WIDTH 11
`define ACC_INT_WIDTH 5
`define ACC_FRACT_WIDTH 6

`define GYRO_WIDTH 14
`define GYRO_INT_WIDTH 6
`define GYRO_FRACT_WIDTH 8

`define ACC_MAG_SQR_WIDTH 16
`define ACC_MAG_SQR_INT_WIDTH 12
`define ACC_MAG_SQR_FRACT_WIDTH 4

`define Q_MAG_SQR_WIDTH 10
`define Q_MAG_SQR_INT_WIDTH 6
`define Q_MAG_SQR_FRACT_WIDTH 4

`define Q_WIDTH 16
`define Q_INT_WIDTH 2
`define Q_FRACT_WIDTH 14

`define Q_TEMP_WIDTH 50
`define Q_TEMP_INT_WIDTH 18
`define Q_TEMP_FRACT_WIDTH 32

`define Q_HALF_WIDTH 16
`define Q_HALF_INT_WIDTH 2
`define Q_HALF_FRACT_WIDTH 14

`define Q_TWO_WIDTH 17
`define Q_TWO_INT_WIDTH 3
`define Q_TWO_FRACT_WIDTH 14

`define Q_DOT_WIDTH 32
`define Q_DOT_INT_WIDTH 16
`define Q_DOT_FRACT_WIDTH 16

`define JACOBIAN_WIDTH 17
`define JACOBIAN_INT_WIDTH 3
`define JACOBIAN_FRACT_WIDTH 14

`define OBJ_FUNC_WIDTH 35
`define OBJ_FUNC_INT_WIDTH 7
`define OBJ_FUNC_FRACT_WIDTH 28

`define Q_HAT_DOT_WIDTH 16
`define Q_HAT_DOT_INT_WIDTH 8
`define Q_HAT_DOT_FRACT_WIDTH 8

`define Q_HAT_DOT_MAG_SQR_WIDTH 16
`define Q_HAT_DOT_MAG_SQR_INT_WIDTH 8
`define Q_HAT_DOT_MAG_SQR_FRACT_WIDTH 8

