`include "madgwickDefines.vh"

`define NUM_ELEMENTS 1000

parameter logic signed [`ACC_WIDTH-1:0] AX_TEST_VECTOR[`NUM_ELEMENTS] = {
    11'b11110111000,
    11'b11110110100,
    11'b11110101101,
    11'b11110100010,
    11'b11110011001,
    11'b11110010000,
    11'b11110001100,
    11'b11110000111,
    11'b11110000100,
    11'b11110000011,
    11'b11110000001,
    11'b11110000011,
    11'b11110000101,
    11'b11110000111,
    11'b11110000110,
    11'b11110000111,
    11'b11110001000,
    11'b11110001100,
    11'b11110001101,
    11'b11110001101,
    11'b11110001011,
    11'b11110000011,
    11'b11101111101,
    11'b11101110110,
    11'b11101101111,
    11'b11101100011,
    11'b11101011010,
    11'b11101001111,
    11'b11101000100,
    11'b11100110111,
    11'b11100101111,
    11'b11100110001,
    11'b11100110000,
    11'b11101001000,
    11'b11101100001,
    11'b11101011000,
    11'b11100100101,
    11'b11011110110,
    11'b11011001010,
    11'b11010101011,
    11'b11010101000,
    11'b11010111001,
    11'b11011001100,
    11'b11011011000,
    11'b11011100010,
    11'b11011100011,
    11'b11011100101,
    11'b11011100111,
    11'b11011101001,
    11'b11011101001,
    11'b11011101000,
    11'b11011101010,
    11'b11011101001,
    11'b11011101010,
    11'b11011101000,
    11'b11011101000,
    11'b11011100111,
    11'b11011100110,
    11'b11011100110,
    11'b11011100001,
    11'b11011011111,
    11'b11011011010,
    11'b11011011010,
    11'b11011010011,
    11'b11011000001,
    11'b11010101100,
    11'b11010100110,
    11'b11010110000,
    11'b11010111011,
    11'b11011001011,
    11'b11011011100,
    11'b11011110111,
    11'b11100001000,
    11'b11100010101,
    11'b11100010111,
    11'b11011101100,
    11'b11010100001,
    11'b11001110100,
    11'b11001011100,
    11'b11001010100,
    11'b11010000100,
    11'b11011101011,
    11'b11101101101,
    11'b11111010100,
    11'b00000001011,
    11'b11110100110,
    11'b11100100010,
    11'b11010111101,
    11'b11010000011,
    11'b11001110110,
    11'b11010010001,
    11'b11010110101,
    11'b11011010011,
    11'b11011100100,
    11'b11011100100,
    11'b11011010100,
    11'b11010111010,
    11'b11010000111,
    11'b11001011010,
    11'b11000110001,
    11'b11000100011,
    11'b11000101010,
    11'b11000011011,
    11'b11000100101,
    11'b11000111101,
    11'b11001011111,
    11'b11011000010,
    11'b11011111100,
    11'b11100100010,
    11'b11101000100,
    11'b11101001011,
    11'b11100011011,
    11'b11011101010,
    11'b11011000110,
    11'b11010111100,
    11'b11011000000,
    11'b11011000110,
    11'b11011000110,
    11'b11011000110,
    11'b11011000100,
    11'b11011000100,
    11'b11010111100,
    11'b11010111101,
    11'b11011000100,
    11'b11011000110,
    11'b11011010101,
    11'b11011011111,
    11'b11011100101,
    11'b11011101100,
    11'b11011110100,
    11'b11011111101,
    11'b11100000100,
    11'b11100010000,
    11'b11100010101,
    11'b11100011101,
    11'b11100011011,
    11'b11100000100,
    11'b11011011011,
    11'b11011001000,
    11'b11011010011,
    11'b11011011000,
    11'b11011010101,
    11'b11011010011,
    11'b11011010100,
    11'b11011000100,
    11'b11011010100,
    11'b11010101011,
    11'b11001100001,
    11'b11010111000,
    11'b11100000110,
    11'b11100000100,
    11'b11011111010,
    11'b11100101101,
    11'b11011100101,
    11'b11011101001,
    11'b11010110011,
    11'b11010010010,
    11'b11010011011,
    11'b11010110110,
    11'b11011001101,
    11'b11011011100,
    11'b11011100000,
    11'b11011010110,
    11'b11011001101,
    11'b11011001110,
    11'b11011100011,
    11'b11011111010,
    11'b11011101100,
    11'b11010111100,
    11'b11010100010,
    11'b11010011000,
    11'b11010011111,
    11'b11010101100,
    11'b11010110010,
    11'b11010110111,
    11'b11011000111,
    11'b11100001001,
    11'b11011111000,
    11'b11011011010,
    11'b11010110011,
    11'b11010111010,
    11'b11011001111,
    11'b11011001010,
    11'b11011111101,
    11'b11100110110,
    11'b11101000011,
    11'b11100001101,
    11'b11011001010,
    11'b11010100011,
    11'b11010101000,
    11'b11011000001,
    11'b11011100011,
    11'b11100001010,
    11'b11100010100,
    11'b11011111111,
    11'b11011011100,
    11'b11010101111,
    11'b11010011100,
    11'b11010010011,
    11'b11010001111,
    11'b11010011010,
    11'b11010111010,
    11'b11010110110,
    11'b11010101001,
    11'b11010111100,
    11'b11010111111,
    11'b11010110101,
    11'b11010111100,
    11'b11011011010,
    11'b11011101010,
    11'b11011101111,
    11'b11011100100,
    11'b11011001111,
    11'b11010110001,
    11'b11010011011,
    11'b11010001010,
    11'b11001111001,
    11'b11001100100,
    11'b11001010001,
    11'b11000111100,
    11'b11000101010,
    11'b11000100001,
    11'b11000101010,
    11'b11000111111,
    11'b11001011100,
    11'b11001110110,
    11'b11010010101,
    11'b11010100010,
    11'b11010101000,
    11'b11010100111,
    11'b11010100011,
    11'b11010100001,
    11'b11010100001,
    11'b11010100011,
    11'b11010100000,
    11'b11010011000,
    11'b11010001010,
    11'b11001111000,
    11'b11001101010,
    11'b11001100001,
    11'b11001011101,
    11'b11001011100,
    11'b11001011100,
    11'b11001011000,
    11'b11001010001,
    11'b11000100110,
    11'b10111111111,
    11'b10101010011,
    11'b10001111101,
    11'b10011001100,
    11'b10100110010,
    11'b10101110010,
    11'b10110100001,
    11'b10111101001,
    11'b11001000011,
    11'b11001100000,
    11'b11010001000,
    11'b11010101000,
    11'b11011010110,
    11'b11011110001,
    11'b11100000011,
    11'b11011111010,
    11'b11011100010,
    11'b11011001111,
    11'b11010110001,
    11'b11010010100,
    11'b11001111000,
    11'b11001100011,
    11'b11001001111,
    11'b11001000100,
    11'b11000111000,
    11'b11000111010,
    11'b11001000100,
    11'b11001010111,
    11'b11001101111,
    11'b11010010100,
    11'b11010101111,
    11'b11010111111,
    11'b11011010111,
    11'b11011110001,
    11'b11100000011,
    11'b11100010100,
    11'b11100010001,
    11'b11011101100,
    11'b11011010110,
    11'b11011001000,
    11'b11010111000,
    11'b11010100000,
    11'b11010001101,
    11'b11010001000,
    11'b11010000110,
    11'b11010001000,
    11'b11010001100,
    11'b11010000100,
    11'b11010000011,
    11'b11010000011,
    11'b11010000110,
    11'b11010001000,
    11'b11010001010,
    11'b11010001010,
    11'b11010001100,
    11'b11010001100,
    11'b11010001101,
    11'b11010010000,
    11'b11010010010,
    11'b11010010100,
    11'b11010010100,
    11'b11010010101,
    11'b11010010011,
    11'b11010010010,
    11'b11010010001,
    11'b11010010000,
    11'b11010001111,
    11'b11010001101,
    11'b11010001100,
    11'b11010001010,
    11'b11010001001,
    11'b11010001000,
    11'b11010001000,
    11'b11010001000,
    11'b11010001000,
    11'b11010001001,
    11'b11010001000,
    11'b11010001011,
    11'b11010001100,
    11'b11010001111,
    11'b11010010000,
    11'b11010010010,
    11'b11010010010,
    11'b11010010011,
    11'b11010010001,
    11'b11010010001,
    11'b11010010001,
    11'b11010010001,
    11'b11010010000,
    11'b11010001111,
    11'b11010001111,
    11'b11010001101,
    11'b11010001101,
    11'b11010001101,
    11'b11010001101,
    11'b11010001101,
    11'b11010001100,
    11'b11010001101,
    11'b11010001100,
    11'b11010001101,
    11'b11010001101,
    11'b11010001110,
    11'b11010001111,
    11'b11010001111,
    11'b11010010000,
    11'b11010010001,
    11'b11010010010,
    11'b11010010001,
    11'b11010010010,
    11'b11010010010,
    11'b11010010011,
    11'b11010010001,
    11'b11010010001,
    11'b11010010001,
    11'b11010001111,
    11'b11010001111,
    11'b11010001111,
    11'b11010001111,
    11'b11010001111,
    11'b11010101000,
    11'b11010111110,
    11'b11011000001,
    11'b11010100100,
    11'b11010011100,
    11'b11010011011,
    11'b11010011000,
    11'b11010011010,
    11'b11010010001,
    11'b11010000100,
    11'b11001110110,
    11'b11001011100,
    11'b11001011101,
    11'b11001100001,
    11'b11001101010,
    11'b11010001000,
    11'b11010010001,
    11'b11010010011,
    11'b11010001111,
    11'b11010000110,
    11'b11010000100,
    11'b11010000100,
    11'b11010001010,
    11'b11010010011,
    11'b11010011001,
    11'b11010011100,
    11'b11010011010,
    11'b11010010110,
    11'b11010010001,
    11'b11010010100,
    11'b11010010111,
    11'b11010011001,
    11'b11010010111,
    11'b11010010011,
    11'b11010010000,
    11'b11010001011,
    11'b11010001011,
    11'b11010001011,
    11'b11010001101,
    11'b11010010000,
    11'b10111100110,
    11'b10111010001,
    11'b11001000100,
    11'b11011011101,
    11'b11001011010,
    11'b11001011100,
    11'b10111101100,
    11'b10110111111,
    11'b10111011100,
    11'b11000000001,
    11'b11000100111,
    11'b11001000011,
    11'b11001100011,
    11'b11001110110,
    11'b11001110101,
    11'b11001110011,
    11'b11001110110,
    11'b11010001100,
    11'b11010110000,
    11'b11000111101,
    11'b11100101101,
    11'b00001001010,
    11'b00010001110,
    11'b00010010001,
    11'b00010001101,
    11'b00010000100,
    11'b00001011000,
    11'b11111011001,
    11'b11100111001,
    11'b11010101001,
    11'b10111110011,
    11'b10101000011,
    11'b10011010010,
    11'b10001111110,
    11'b10000111111,
    11'b10000101000,
    11'b10001000011,
    11'b10001100100,
    11'b10010100001,
    11'b10100000100,
    11'b10101100100,
    11'b10111001010,
    11'b11001011011,
    11'b11010101100,
    11'b11011110001,
    11'b11100100011,
    11'b11101010111,
    11'b11101111010,
    11'b11110011000,
    11'b11110110100,
    11'b11111000101,
    11'b11110111100,
    11'b11110000001,
    11'b11101100001,
    11'b11100111010,
    11'b11100000001,
    11'b11011110000,
    11'b11011100011,
    11'b11011001100,
    11'b11010100011,
    11'b11010000011,
    11'b11001100100,
    11'b11001011100,
    11'b11001101000,
    11'b11001110000,
    11'b11001110101,
    11'b11001111000,
    11'b11001110010,
    11'b11001101010,
    11'b11001100100,
    11'b11001011101,
    11'b11010001000,
    11'b11010011010,
    11'b11010011101,
    11'b11010100000,
    11'b11010011000,
    11'b11010000100,
    11'b11001111110,
    11'b11010000000,
    11'b11010001001,
    11'b11010010100,
    11'b11010010011,
    11'b11010010001,
    11'b11010001111,
    11'b11010001000,
    11'b11010001000,
    11'b11010001000,
    11'b11010010000,
    11'b11010010110,
    11'b11010011100,
    11'b11010100001,
    11'b11010100011,
    11'b11010100111,
    11'b11010100111,
    11'b11010101010,
    11'b11010101010,
    11'b11010101011,
    11'b11010101001,
    11'b11010100011,
    11'b11010011101,
    11'b11010010110,
    11'b11010010001,
    11'b11010011010,
    11'b11010011110,
    11'b11010001010,
    11'b11001111111,
    11'b11010000001,
    11'b11001101001,
    11'b11001100111,
    11'b11001101100,
    11'b11100111111,
    11'b00100000110,
    11'b00000010011,
    11'b11010010011,
    11'b11001011101,
    11'b11000011010,
    11'b11010001000,
    11'b11001001111,
    11'b11000000100,
    11'b10111100110,
    11'b11000111001,
    11'b11010000011,
    11'b11010001001,
    11'b11010101010,
    11'b11010100100,
    11'b11001101010,
    11'b11000110010,
    11'b11000011111,
    11'b11000001101,
    11'b11000100110,
    11'b11001000100,
    11'b11001001111,
    11'b11001111110,
    11'b11011101100,
    11'b11101101000,
    11'b11101110100,
    11'b11011000100,
    11'b11000010000,
    11'b10110000100,
    11'b10101001110,
    11'b10110001100,
    11'b10111100000,
    11'b11000100100,
    11'b11001000001,
    11'b11000111000,
    11'b11000011101,
    11'b11000010000,
    11'b11000010100,
    11'b11000011110,
    11'b11000011101,
    11'b11000010001,
    11'b11000010010,
    11'b11000100001,
    11'b11000101111,
    11'b11000111110,
    11'b11001001000,
    11'b11001001101,
    11'b11001001101,
    11'b11001001000,
    11'b11001001011,
    11'b11001010100,
    11'b11001011000,
    11'b11001010100,
    11'b11001010001,
    11'b11001001101,
    11'b11000111111,
    11'b11000100011,
    11'b11000000001,
    11'b10111101000,
    11'b10111011010,
    11'b10111010010,
    11'b10111001010,
    11'b10111000000,
    11'b10110111101,
    11'b10111000001,
    11'b10111001000,
    11'b10111011000,
    11'b10111101001,
    11'b10111111001,
    11'b11000001000,
    11'b11000010100,
    11'b11000110110,
    11'b11001001001,
    11'b11001010110,
    11'b11001100011,
    11'b11001110100,
    11'b11001000100,
    11'b11000100100,
    11'b11000111111,
    11'b11010000001,
    11'b11010111010,
    11'b11011100100,
    11'b11011111010,
    11'b11100000100,
    11'b11100000111,
    11'b11100011011,
    11'b11100101000,
    11'b11100110001,
    11'b11101001011,
    11'b11101010111,
    11'b11101001000,
    11'b11101010110,
    11'b11101010110,
    11'b11101011011,
    11'b11101100100,
    11'b11101011111,
    11'b11101010110,
    11'b11101010010,
    11'b11101000100,
    11'b11101001010,
    11'b11101001000,
    11'b11101001111,
    11'b11101000001,
    11'b11101000001,
    11'b11100111111,
    11'b11100100000,
    11'b11100011010,
    11'b11100101101,
    11'b11100111011,
    11'b11101010010,
    11'b11100101011,
    11'b11100001100,
    11'b11011110100,
    11'b11100011010,
    11'b00001000100,
    11'b00111100100,
    11'b01001111010,
    11'b00110111000,
    11'b00100100111,
    11'b00011010110,
    11'b00010011000,
    11'b00000011111,
    11'b00000000001,
    11'b00001001101,
    11'b00010111011,
    11'b00100000010,
    11'b00100101000,
    11'b00100111111,
    11'b00101000000,
    11'b00100011111,
    11'b00011101100,
    11'b00011011100,
    11'b00011010000,
    11'b00010111010,
    11'b00010011001,
    11'b00010001101,
    11'b00010010001,
    11'b00010010011,
    11'b00010010001,
    11'b00010011001,
    11'b00001111111,
    11'b00001001101,
    11'b11111110100,
    11'b11110001111,
    11'b11101110111,
    11'b11110100011,
    11'b11111010001,
    11'b00000001111,
    11'b00001011100,
    11'b00001110000,
    11'b00001110100,
    11'b00010000001,
    11'b00010010011,
    11'b00010100001,
    11'b00010100010,
    11'b00010001010,
    11'b00001110010,
    11'b00001110001,
    11'b00010000100,
    11'b00010010110,
    11'b00010100100,
    11'b00010101111,
    11'b00010110011,
    11'b00010110001,
    11'b00010100011,
    11'b00010100110,
    11'b00011000111,
    11'b00100010001,
    11'b00101011111,
    11'b00110001010,
    11'b00110111001,
    11'b00111001000,
    11'b00111011101,
    11'b00111100101,
    11'b00111000100,
    11'b00110011100,
    11'b00101110011,
    11'b00101000110,
    11'b00100000001,
    11'b00011101111,
    11'b00011111011,
    11'b00100010111,
    11'b00100110100,
    11'b00101000001,
    11'b00101000110,
    11'b00101001101,
    11'b00101010100,
    11'b00101010110,
    11'b00101001111,
    11'b00101000001,
    11'b00100110010,
    11'b00100011010,
    11'b00100001001,
    11'b00011111000,
    11'b00011101000,
    11'b00011100110,
    11'b00011101100,
    11'b00011110100,
    11'b00011110110,
    11'b00011110110,
    11'b00011110011,
    11'b00011111111,
    11'b00011101111,
    11'b00011111010,
    11'b00011111000,
    11'b00100001010,
    11'b00100011001,
    11'b00100011101,
    11'b00100001100,
    11'b00100010100,
    11'b00100001000,
    11'b00100000101,
    11'b00100001101,
    11'b00100000001,
    11'b00011100011,
    11'b00011000111,
    11'b00010100111,
    11'b00100111001,
    11'b00010101001,
    11'b00000100000,
    11'b00000110001,
    11'b00001011001,
    11'b00000001011,
    11'b11111010110,
    11'b00000111001,
    11'b00010110001,
    11'b00010010101,
    11'b00001101000,
    11'b00000111110,
    11'b00000011010,
    11'b11111111101,
    11'b11111111111,
    11'b00000001001,
    11'b00000010100,
    11'b00000010100,
    11'b00000011000,
    11'b00000011101,
    11'b00000100100,
    11'b00000101011,
    11'b00000110001,
    11'b00000110100,
    11'b00000111000,
    11'b00001001111,
    11'b00001011101,
    11'b00001101000,
    11'b00001111111,
    11'b00010011000,
    11'b00010100000,
    11'b00010101010,
    11'b00011001000,
    11'b00011001100,
    11'b00011011111,
    11'b00011100010,
    11'b00011110100,
    11'b00011110110,
    11'b00011111100,
    11'b00100000000,
    11'b00011111111,
    11'b00011111110,
    11'b00011111001,
    11'b00011111111,
    11'b00011111110,
    11'b00011110011,
    11'b00011011000,
    11'b00010101111,
    11'b00010010001,
    11'b00001101101,
    11'b00001001101,
    11'b00000111110,
    11'b00000101001,
    11'b00000101111,
    11'b00000100110,
    11'b00000010101,
    11'b00000110101,
    11'b00001011101,
    11'b00001101010,
    11'b00001101000,
    11'b00001110001,
    11'b00010000001,
    11'b00010010001,
    11'b00010011000,
    11'b00010100011,
    11'b00010110001,
    11'b00010111111,
    11'b00011001100,
    11'b00011010011,
    11'b00011100010,
    11'b00011101101,
    11'b00011111010,
    11'b00100001000,
    11'b00100011001,
    11'b00100100101,
    11'b00100101110,
    11'b00100101111,
    11'b00100110011,
    11'b00100110000,
    11'b00100100100,
    11'b00100010110,
    11'b00100001100,
    11'b00011100110,
    11'b00011101110,
    11'b00011011111,
    11'b00011000100,
    11'b00010110011,
    11'b00011001110,
    11'b00010100000,
    11'b00010110000,
    11'b00011000000,
    11'b00010111011,
    11'b00010110011,
    11'b00010101010,
    11'b00010100011,
    11'b00010010100,
    11'b00010001101,
    11'b00010001111,
    11'b00010001100,
    11'b00010001100,
    11'b00010000110,
    11'b00001111111,
    11'b00001110101,
    11'b00001111000,
    11'b00001101111,
    11'b00001101001,
    11'b00001100011,
    11'b00001100001,
    11'b00001011010,
    11'b00001010101,
    11'b00001001000,
    11'b00000111101,
    11'b00000110101,
    11'b00000100011,
    11'b00000011101,
    11'b00000011000,
    11'b00000010010,
    11'b00000001101,
    11'b00000001100,
    11'b00000001100,
    11'b00000001011,
    11'b00000001110,
    11'b00000010001,
    11'b00000010011,
    11'b00000010110,
    11'b00000011101,
    11'b00000011111,
    11'b00000100000,
    11'b00000011110,
    11'b00000010111,
    11'b00000010011,
    11'b00000001110,
    11'b00000001000,
    11'b00000000001,
    11'b11111111000,
    11'b11111110001,
    11'b11111101011,
    11'b11111101000,
    11'b11111100100,
    11'b11111100011,
    11'b11111100000,
    11'b11111100001,
    11'b11111100000,
    11'b11111100111,
    11'b11111110011,
    11'b11111111100,
    11'b00000000001,
    11'b00000000011,
    11'b00000001000,
    11'b00000010001,
    11'b00000001100,
    11'b11111111111,
    11'b11111110110,
    11'b11111110110,
    11'b11111110011,
    11'b11111101010,
    11'b11111100101,
    11'b11111011001,
    11'b11111011100,
    11'b11111010110,
    11'b11111010011,
    11'b11111000110,
    11'b11110111010,
    11'b11110010100,
    11'b11110100110,
    11'b11110101011,
    11'b11110100100,
    11'b11110101100,
    11'b11110110011,
    11'b11110111100,
    11'b11110110010,
    11'b11110111001,
    11'b11111011000,
    11'b11111011011,
    11'b11111010110,
    11'b11111000001,
    11'b11101001001,
    11'b11011001101,
    11'b11010001001,
    11'b11001111000,
    11'b10111100101,
    11'b10110001101,
    11'b10111100110,
    11'b11010011100,
    11'b11100110110,
    11'b11110101111,
    11'b00110001100,
    11'b01010100100,
    11'b01101000010,
    11'b01011010001,
    11'b00111001000,
    11'b00100010110,
    11'b00010011101,
    11'b00000101111,
    11'b11110011101,
    11'b11101101101,
    11'b11101111100,
    11'b11110101001,
    11'b11110001101,
    11'b11101011111,
    11'b11101000000,
    11'b11101110100,
    11'b11111110111,
    11'b00000011000,
    11'b00000100001,
    11'b00000100011,
    11'b00000100000,
    11'b00010001101,
    11'b00010010110,
    11'b00001001010,
    11'b11111101111,
    11'b11111001111,
    11'b11110111001,
    11'b11111000100,
    11'b11111011101,
    11'b11111111101,
    11'b11110111000,
    11'b11101100111,
    11'b11110000010,
    11'b11101111010,
    11'b11101100110,
    11'b11101011011,
    11'b11101101110,
    11'b11110101001,
    11'b11110101100,
    11'b11101100100,
    11'b11101111100,
    11'b11110100101,
    11'b11110110110,
    11'b11111001000,
    11'b11111110001,
    11'b00001000110,
    11'b00011000110,
    11'b00101110101,
    11'b00110100001,
    11'b00101010100,
    11'b00100000110,
    11'b00011111000,
    11'b00100111101,
    11'b00100100001,
    11'b00100011010,
    11'b00011011000,
    11'b00101011000,
    11'b00100101100,
    11'b01010000100,
    11'b00111110100,
    11'b00110010110,
    11'b00101111111,
    11'b00101100011,
    11'b00110000001,
    11'b00110011111,
    11'b00110001011,
    11'b00110001000,
    11'b00101100011,
    11'b00101000110,
    11'b00100110110,
    11'b00100110110,
    11'b00100110011,
    11'b00100111000,
    11'b00100111001,
    11'b00100110011,
    11'b00101000101,
    11'b00101010100,
    11'b00110100001,
    11'b00111010011,
    11'b01000001110,
    11'b01001001100,
    11'b01010000110
};

parameter logic signed [`ACC_WIDTH-1:0] AY_TEST_VECTOR[`NUM_ELEMENTS] = {
    11'b00101001010,
    11'b00101001001,
    11'b00101000110,
    11'b00101000001,
    11'b00100111101,
    11'b00100110110,
    11'b00100110010,
    11'b00100101110,
    11'b00100101010,
    11'b00100011111,
    11'b00100010101,
    11'b00100001110,
    11'b00100001100,
    11'b00100001100,
    11'b00100001010,
    11'b00100001001,
    11'b00100000100,
    11'b00011111111,
    11'b00011111010,
    11'b00011110100,
    11'b00011110000,
    11'b00011101000,
    11'b00011100010,
    11'b00011011101,
    11'b00011011001,
    11'b00011010011,
    11'b00011001101,
    11'b00011001000,
    11'b00011000001,
    11'b00010110101,
    11'b00010101010,
    11'b00010011110,
    11'b00010001110,
    11'b00010000001,
    11'b00001110111,
    11'b00001101010,
    11'b00001010110,
    11'b00001001111,
    11'b00001001101,
    11'b00001010001,
    11'b00001010011,
    11'b00001001101,
    11'b00001000011,
    11'b00000110111,
    11'b00000101111,
    11'b00000101010,
    11'b00000101000,
    11'b00000100100,
    11'b00000011100,
    11'b00000010011,
    11'b00000001011,
    11'b00000000110,
    11'b11111111111,
    11'b11111111010,
    11'b11111110110,
    11'b11111110001,
    11'b11111101110,
    11'b11111101101,
    11'b11111101100,
    11'b11111101101,
    11'b11111101111,
    11'b11111110000,
    11'b11111110010,
    11'b11111110010,
    11'b11111100011,
    11'b11111010100,
    11'b11111010001,
    11'b11111011000,
    11'b11111011100,
    11'b11111100100,
    11'b11111110000,
    11'b11111111101,
    11'b00000001011,
    11'b00000010100,
    11'b00000100000,
    11'b00001001101,
    11'b00010010000,
    11'b00010110001,
    11'b00011011101,
    11'b00100001101,
    11'b00100110101,
    11'b00011110010,
    11'b00001100110,
    11'b11111001101,
    11'b11101100101,
    11'b11101011000,
    11'b11110100011,
    11'b11111110001,
    11'b00000010110,
    11'b00000011001,
    11'b00000010111,
    11'b00000100001,
    11'b00000110001,
    11'b00000111010,
    11'b00000101010,
    11'b00000001110,
    11'b11111101111,
    11'b11111011010,
    11'b11111100000,
    11'b11111101001,
    11'b11111101011,
    11'b11111110110,
    11'b00000000111,
    11'b00000100011,
    11'b00000111100,
    11'b00001010011,
    11'b00001111000,
    11'b00010001000,
    11'b00010001111,
    11'b00010011001,
    11'b00010011000,
    11'b00010000001,
    11'b00001101000,
    11'b00001011011,
    11'b00001011011,
    11'b00001100011,
    11'b00001100111,
    11'b00001101001,
    11'b00001101011,
    11'b00001101101,
    11'b00001101110,
    11'b00010001111,
    11'b00010110010,
    11'b00010000110,
    11'b00001011101,
    11'b00001011110,
    11'b00001010110,
    11'b00001010110,
    11'b00001101000,
    11'b00001101110,
    11'b00001110000,
    11'b00001101111,
    11'b00001100011,
    11'b00001100011,
    11'b00001100000,
    11'b00001011001,
    11'b00001100001,
    11'b00001101110,
    11'b00001100100,
    11'b00001011110,
    11'b00000111110,
    11'b00000100011,
    11'b00000001011,
    11'b00000001011,
    11'b00000001101,
    11'b00000010011,
    11'b00000011000,
    11'b00000011110,
    11'b00001000001,
    11'b00001001100,
    11'b00001010000,
    11'b00001010001,
    11'b00000111110,
    11'b00000110011,
    11'b00000101100,
    11'b00000101000,
    11'b00000111101,
    11'b00001011100,
    11'b00001111100,
    11'b00010010001,
    11'b00010010110,
    11'b00010001100,
    11'b00010000001,
    11'b00001111010,
    11'b00001101011,
    11'b00001100100,
    11'b00001011010,
    11'b00001100101,
    11'b00001101101,
    11'b00001010110,
    11'b00000111000,
    11'b00000100010,
    11'b00000010010,
    11'b00000000110,
    11'b11111111000,
    11'b11111101001,
    11'b11111010111,
    11'b11111010110,
    11'b11111100100,
    11'b11111010001,
    11'b11110101110,
    11'b11110100110,
    11'b11111001100,
    11'b00000010101,
    11'b00001010100,
    11'b00010010111,
    11'b00011010100,
    11'b00100000100,
    11'b00100100110,
    11'b00100100010,
    11'b00100011000,
    11'b00100010100,
    11'b00100001001,
    11'b00011110011,
    11'b00011001001,
    11'b00010001111,
    11'b00000110010,
    11'b11111101101,
    11'b11110101011,
    11'b11101110100,
    11'b11100110001,
    11'b11011110110,
    11'b11011100110,
    11'b11011100101,
    11'b11011001111,
    11'b11010111101,
    11'b11011001000,
    11'b11011001100,
    11'b11011100101,
    11'b11100000111,
    11'b11100101010,
    11'b11101001010,
    11'b11101100111,
    11'b11110000010,
    11'b11110001111,
    11'b11110011000,
    11'b11110100000,
    11'b11110110011,
    11'b11111001000,
    11'b11111100010,
    11'b11111111101,
    11'b00000011110,
    11'b00000101110,
    11'b00000110010,
    11'b00000101010,
    11'b00000010111,
    11'b11111111000,
    11'b11111100010,
    11'b11111010001,
    11'b11111000110,
    11'b11111000011,
    11'b11111000110,
    11'b11111001100,
    11'b11111010011,
    11'b11111011010,
    11'b11111100001,
    11'b11111100110,
    11'b11111101101,
    11'b11111110010,
    11'b11111111000,
    11'b11111111111,
    11'b00000010001,
    11'b00000100100,
    11'b00000111011,
    11'b00001010000,
    11'b00001010111,
    11'b00001000111,
    11'b00000101111,
    11'b11111100110,
    11'b00000101101,
    11'b00000111011,
    11'b00001011100,
    11'b00001001011,
    11'b00001011000,
    11'b00001000100,
    11'b00001011010,
    11'b00001101100,
    11'b00001011010,
    11'b00000010010,
    11'b11111010101,
    11'b11110000100,
    11'b11101000110,
    11'b11100010111,
    11'b11100011101,
    11'b11100111010,
    11'b11101010001,
    11'b11101011011,
    11'b11101010101,
    11'b11101000111,
    11'b11100111000,
    11'b11100101110,
    11'b11100010110,
    11'b11100001011,
    11'b11100001000,
    11'b11100001111,
    11'b11100010110,
    11'b11100100011,
    11'b11100110010,
    11'b11100111000,
    11'b11100111111,
    11'b11101000011,
    11'b11101001001,
    11'b11101001111,
    11'b11101100100,
    11'b11110001100,
    11'b11110101010,
    11'b11110111101,
    11'b11111010100,
    11'b11111011101,
    11'b11111100011,
    11'b11111100110,
    11'b11111101000,
    11'b11111101000,
    11'b11111101011,
    11'b11111101011,
    11'b11111101010,
    11'b11111101010,
    11'b11111101010,
    11'b11111101010,
    11'b11111101001,
    11'b11111101010,
    11'b11111101010,
    11'b11111101010,
    11'b11111101010,
    11'b11111101010,
    11'b11111101011,
    11'b11111101100,
    11'b11111101100,
    11'b11111101100,
    11'b11111101101,
    11'b11111101100,
    11'b11111101100,
    11'b11111101100,
    11'b11111101100,
    11'b11111101101,
    11'b11111101101,
    11'b11111101100,
    11'b11111101100,
    11'b11111101101,
    11'b11111101100,
    11'b11111101011,
    11'b11111101011,
    11'b11111101011,
    11'b11111101011,
    11'b11111101010,
    11'b11111101011,
    11'b11111101010,
    11'b11111101010,
    11'b11111101011,
    11'b11111101011,
    11'b11111101011,
    11'b11111101100,
    11'b11111101010,
    11'b11111101011,
    11'b11111101011,
    11'b11111101010,
    11'b11111101011,
    11'b11111101010,
    11'b11111101100,
    11'b11111101100,
    11'b11111101011,
    11'b11111101010,
    11'b11111101010,
    11'b11111101010,
    11'b11111101010,
    11'b11111101010,
    11'b11111101000,
    11'b11111101000,
    11'b11111101001,
    11'b11111101010,
    11'b11111101010,
    11'b11111101001,
    11'b11111101001,
    11'b11111101000,
    11'b11111101000,
    11'b11111101001,
    11'b11111101001,
    11'b11111101001,
    11'b11111101010,
    11'b11111101010,
    11'b11111101010,
    11'b11111101010,
    11'b11111101010,
    11'b11111101010,
    11'b11111101010,
    11'b11111101110,
    11'b11111110011,
    11'b11111110100,
    11'b11111110001,
    11'b11111110011,
    11'b11111111010,
    11'b00000000011,
    11'b00000001001,
    11'b00000000101,
    11'b11111110011,
    11'b11111011100,
    11'b11111000100,
    11'b11111001111,
    11'b11111010110,
    11'b11111011111,
    11'b11111100110,
    11'b11111101000,
    11'b11111100111,
    11'b11111101010,
    11'b11111101000,
    11'b11111101001,
    11'b11111101010,
    11'b11111101010,
    11'b11111101000,
    11'b11111101010,
    11'b11111101010,
    11'b11111101010,
    11'b11111101100,
    11'b11111101010,
    11'b11111101011,
    11'b11111101011,
    11'b11111101100,
    11'b11111101100,
    11'b11111101011,
    11'b11111101010,
    11'b11111101001,
    11'b11111101001,
    11'b11111101010,
    11'b11111101001,
    11'b11111101001,
    11'b10000000000,
    11'b10000000000,
    11'b10110000111,
    11'b01111100011,
    11'b00110111000,
    11'b00100010011,
    11'b00010010101,
    11'b00000100111,
    11'b11111110111,
    11'b11111011101,
    11'b11111010011,
    11'b11110111111,
    11'b11111000010,
    11'b11110100110,
    11'b11111010001,
    11'b11111111000,
    11'b00000111001,
    11'b00010100110,
    11'b00110010110,
    11'b01011000111,
    11'b01011011000,
    11'b01011001001,
    11'b01001011010,
    11'b01000000001,
    11'b00110110100,
    11'b00110000111,
    11'b00100111110,
    11'b00010101010,
    11'b00001100001,
    11'b00000000010,
    11'b11110001010,
    11'b11010110100,
    11'b11001101110,
    11'b11000111011,
    11'b11000011001,
    11'b11000001010,
    11'b11000010011,
    11'b11000110001,
    11'b11001011000,
    11'b11010010111,
    11'b11011010011,
    11'b11100010010,
    11'b11101110001,
    11'b11110101010,
    11'b11111010101,
    11'b11111110110,
    11'b00000001101,
    11'b00000011101,
    11'b00000101011,
    11'b00000110011,
    11'b00000100111,
    11'b00000000010,
    11'b11111010111,
    11'b11111001010,
    11'b11110111101,
    11'b11111000100,
    11'b11111011100,
    11'b11111101011,
    11'b11111101100,
    11'b11111100011,
    11'b11111011000,
    11'b11111010011,
    11'b11111011001,
    11'b11111110001,
    11'b00000000000,
    11'b00000001100,
    11'b00000010001,
    11'b00000010001,
    11'b00000001011,
    11'b00000001001,
    11'b11111111111,
    11'b11111101101,
    11'b11111100110,
    11'b11111100100,
    11'b11111100011,
    11'b11111101101,
    11'b11111101000,
    11'b11111100110,
    11'b11111110110,
    11'b00000000111,
    11'b00000000110,
    11'b00000000010,
    11'b11111111101,
    11'b11111111010,
    11'b11111110111,
    11'b11111110110,
    11'b11111110110,
    11'b11111111001,
    11'b11111111000,
    11'b11111110110,
    11'b11111110110,
    11'b11111110011,
    11'b11111110001,
    11'b11111101110,
    11'b11111101100,
    11'b11111101010,
    11'b11111101000,
    11'b11111101001,
    11'b11111110001,
    11'b11111111000,
    11'b11111110100,
    11'b11111110100,
    11'b11111110100,
    11'b11111110100,
    11'b11111111111,
    11'b00000010011,
    11'b00000011100,
    11'b00000100000,
    11'b00000011111,
    11'b00000011101,
    11'b11101001000,
    11'b10001010111,
    11'b10001100000,
    11'b11000000111,
    11'b11010001011,
    11'b11100001111,
    11'b00011011101,
    11'b00010101101,
    11'b00001110001,
    11'b00000110100,
    11'b11111011100,
    11'b11110001010,
    11'b11100111100,
    11'b11100111000,
    11'b11100110001,
    11'b11100100100,
    11'b11100011001,
    11'b11100101101,
    11'b11101101111,
    11'b11110101101,
    11'b11111001101,
    11'b11111101100,
    11'b00100111111,
    11'b01100010001,
    11'b01111111111,
    11'b01111111111,
    11'b01011110001,
    11'b00101000001,
    11'b11111100100,
    11'b11100011100,
    11'b11100000100,
    11'b11101111111,
    11'b00000101110,
    11'b00010111110,
    11'b00011110111,
    11'b00010111111,
    11'b00001111000,
    11'b00001011100,
    11'b00001111111,
    11'b00011001001,
    11'b00011010011,
    11'b00011101110,
    11'b00100011111,
    11'b00100111100,
    11'b00100110111,
    11'b00100011101,
    11'b00100000110,
    11'b00011111100,
    11'b00100000000,
    11'b00100001111,
    11'b00100100010,
    11'b00100011111,
    11'b00100101011,
    11'b00100111000,
    11'b00100101101,
    11'b00100011100,
    11'b00011111100,
    11'b00011001000,
    11'b00010101011,
    11'b00010001010,
    11'b00001110100,
    11'b00001100110,
    11'b00001010101,
    11'b00001001010,
    11'b00001001100,
    11'b00001011001,
    11'b00001100001,
    11'b00001100011,
    11'b00001011001,
    11'b00001010000,
    11'b00001001100,
    11'b00001001110,
    11'b00001011010,
    11'b00001100000,
    11'b00001110100,
    11'b00001111000,
    11'b11110010111,
    11'b11011000001,
    11'b11010101101,
    11'b11110011000,
    11'b00010001001,
    11'b00101101101,
    11'b00111111111,
    11'b01000011110,
    11'b01000011010,
    11'b01000110001,
    11'b01000101101,
    11'b01000000100,
    11'b01000010101,
    11'b00111101000,
    11'b00110011100,
    11'b00110001101,
    11'b00100001000,
    11'b00101011000,
    11'b00110101000,
    11'b00110101111,
    11'b00110011011,
    11'b00100100011,
    11'b00011010111,
    11'b00001110001,
    11'b00000101111,
    11'b11111011010,
    11'b11110111000,
    11'b11110101010,
    11'b11110100110,
    11'b11110010011,
    11'b11101111111,
    11'b11101110011,
    11'b11101001111,
    11'b11100011000,
    11'b11011110111,
    11'b11011101101,
    11'b11011010110,
    11'b11011100011,
    11'b00001011101,
    11'b01010111010,
    11'b01111111111,
    11'b01111111111,
    11'b01111111111,
    11'b01111111111,
    11'b01111110011,
    11'b01011000011,
    11'b00111100001,
    11'b00100101100,
    11'b00010001010,
    11'b00000100100,
    11'b00000100011,
    11'b00001110010,
    11'b00010011111,
    11'b00010001001,
    11'b00001010101,
    11'b00001000100,
    11'b00001000101,
    11'b00001001101,
    11'b00001100100,
    11'b00011000100,
    11'b00100001011,
    11'b00101001001,
    11'b00101101001,
    11'b00110011001,
    11'b00110010111,
    11'b00101101110,
    11'b00100111011,
    11'b00100101000,
    11'b00100011101,
    11'b00100000100,
    11'b00011110100,
    11'b00011111000,
    11'b00100101011,
    11'b00101010001,
    11'b00110000001,
    11'b00110101101,
    11'b00110111101,
    11'b00110010100,
    11'b00101110011,
    11'b00101001101,
    11'b00100110111,
    11'b00100100110,
    11'b00100001110,
    11'b00011101110,
    11'b00011001010,
    11'b00010011101,
    11'b00010000110,
    11'b00001111111,
    11'b00010001010,
    11'b00010011011,
    11'b00011000100,
    11'b00011101111,
    11'b00100101010,
    11'b00101100101,
    11'b00110111111,
    11'b00111110100,
    11'b01000110100,
    11'b01001101110,
    11'b01010110000,
    11'b01011110011,
    11'b01100101100,
    11'b01101010101,
    11'b01101101100,
    11'b01101110000,
    11'b01101101100,
    11'b01101100110,
    11'b01101011000,
    11'b01101000110,
    11'b01100110011,
    11'b01100100101,
    11'b01100101011,
    11'b01100111101,
    11'b01101000011,
    11'b01100111100,
    11'b01100101111,
    11'b01100011100,
    11'b01100010001,
    11'b01100000110,
    11'b01011111101,
    11'b01011110001,
    11'b01011100011,
    11'b01011100000,
    11'b01011100001,
    11'b01011101010,
    11'b01100000011,
    11'b01101000001,
    11'b01101000011,
    11'b01100111101,
    11'b01100110001,
    11'b01100110011,
    11'b01101000001,
    11'b01101100101,
    11'b01101000101,
    11'b01101010001,
    11'b01101101101,
    11'b01101101011,
    11'b01101100100,
    11'b01101101100,
    11'b01101101000,
    11'b01101000111,
    11'b01011011010,
    11'b01001100111,
    11'b01010101011,
    11'b01011110011,
    11'b01011010110,
    11'b01010110100,
    11'b01010100011,
    11'b01001100100,
    11'b01000001000,
    11'b00111000111,
    11'b01000001101,
    11'b01001010000,
    11'b01001111111,
    11'b01010100010,
    11'b01010101010,
    11'b01010100001,
    11'b01010010100,
    11'b01010000110,
    11'b01001111100,
    11'b01001110000,
    11'b01001101111,
    11'b01001011110,
    11'b01001001000,
    11'b01001001010,
    11'b01000110101,
    11'b01000101111,
    11'b01000110001,
    11'b01000111001,
    11'b01000110110,
    11'b01000110011,
    11'b01000111110,
    11'b01000110101,
    11'b01000101010,
    11'b01000110110,
    11'b01000111110,
    11'b01001010011,
    11'b01001000000,
    11'b01000111010,
    11'b01000011010,
    11'b01000000100,
    11'b00111110110,
    11'b00111100000,
    11'b00110111010,
    11'b00110011101,
    11'b00110000011,
    11'b00101101000,
    11'b00101010111,
    11'b00101010101,
    11'b00101010011,
    11'b00101010001,
    11'b00101010100,
    11'b00101001101,
    11'b00101000010,
    11'b00100110110,
    11'b00100011100,
    11'b00100001011,
    11'b00011110001,
    11'b00011011111,
    11'b00011010100,
    11'b00011001101,
    11'b00011000100,
    11'b00010101100,
    11'b00010010100,
    11'b00010000011,
    11'b00001110000,
    11'b00001001100,
    11'b00000101100,
    11'b00000001111,
    11'b11111110110,
    11'b11111100010,
    11'b11111010001,
    11'b11111001000,
    11'b11111000011,
    11'b11110111100,
    11'b11110101100,
    11'b11110011101,
    11'b11110001000,
    11'b11101101111,
    11'b11101001110,
    11'b11100111001,
    11'b11100101011,
    11'b11100100000,
    11'b11100001101,
    11'b11100000111,
    11'b11011011111,
    11'b11010110101,
    11'b11010011101,
    11'b11001101101,
    11'b11001000110,
    11'b11000110000,
    11'b11000000100,
    11'b10111100001,
    11'b10111001000,
    11'b10110110000,
    11'b10110011101,
    11'b10110001110,
    11'b10101111010,
    11'b10101101111,
    11'b10101100101,
    11'b10101100001,
    11'b10101011011,
    11'b10101011100,
    11'b10101011100,
    11'b10101100011,
    11'b10101100110,
    11'b10101101101,
    11'b10101110100,
    11'b10101110101,
    11'b10101110110,
    11'b10101110011,
    11'b10101101111,
    11'b10101101111,
    11'b10101101011,
    11'b10101101001,
    11'b10101100100,
    11'b10101100000,
    11'b10101011101,
    11'b10101011110,
    11'b10101100000,
    11'b10101100101,
    11'b10101101011,
    11'b10101110000,
    11'b10101111001,
    11'b10101111010,
    11'b10101111100,
    11'b10101110111,
    11'b10101101010,
    11'b10101011101,
    11'b10101001111,
    11'b10100111111,
    11'b10100110110,
    11'b10100100101,
    11'b10100011011,
    11'b10100010100,
    11'b10100001111,
    11'b10100001100,
    11'b10100001100,
    11'b10100010010,
    11'b10100011000,
    11'b10100100000,
    11'b10100101110,
    11'b10100111011,
    11'b10101001010,
    11'b10101011100,
    11'b10101111001,
    11'b10110010100,
    11'b10110100111,
    11'b10110111000,
    11'b10111011100,
    11'b10111100010,
    11'b10111001001,
    11'b10111000001,
    11'b10111001001,
    11'b10111001101,
    11'b10110111000,
    11'b10110110001,
    11'b10110111001,
    11'b10110101111,
    11'b10110111001,
    11'b10110110011,
    11'b10110101111,
    11'b10111000111,
    11'b10111011111,
    11'b10111111000,
    11'b11000010010,
    11'b11000100100,
    11'b11000110110,
    11'b11001010010,
    11'b11001110001,
    11'b11010100011,
    11'b11011001100,
    11'b11100010110,
    11'b11110001011,
    11'b11111101010,
    11'b00000001000,
    11'b00000011010,
    11'b00001000100,
    11'b00011101100,
    11'b00101111011,
    11'b00111011100,
    11'b00110100110,
    11'b00000010001,
    11'b11011100111,
    11'b11011010111,
    11'b11101101110,
    11'b00001111100,
    11'b01111111111,
    11'b01010000011,
    11'b00010011101,
    11'b00000010010,
    11'b00000010001,
    11'b11110100001,
    11'b11011101110,
    11'b11011000111,
    11'b11100000001,
    11'b11101110001,
    11'b11110111010,
    11'b11111100110,
    11'b00000000011,
    11'b11110110010,
    11'b11110011111,
    11'b11110100000,
    11'b11110101111,
    11'b11111100011,
    11'b11110100100,
    11'b11110010001,
    11'b11111000011,
    11'b00001011000,
    11'b00011110001,
    11'b00100100101,
    11'b00011011101,
    11'b00010011000,
    11'b00001110011,
    11'b00000100111,
    11'b11111011111,
    11'b11101011000,
    11'b11011000110,
    11'b11001111001,
    11'b11001000001,
    11'b11001010110,
    11'b11010001111,
    11'b11010000110,
    11'b11010000010,
    11'b11011101100,
    11'b11100101111,
    11'b11110100010,
    11'b00000111111,
    11'b00000111111,
    11'b11110011111,
    11'b11100111000,
    11'b11110010110,
    11'b11110110001,
    11'b11110001101,
    11'b11101110000,
    11'b11101010010,
    11'b11101011101,
    11'b11110000110,
    11'b11101111100,
    11'b11101000101,
    11'b11100010100,
    11'b11011011011,
    11'b11011010111,
    11'b11011001110,
    11'b11100001001,
    11'b11011111000,
    11'b11100001000,
    11'b11010111001,
    11'b11011111100,
    11'b11100101111,
    11'b11101101111,
    11'b11111000010,
    11'b11111010100,
    11'b11111001010,
    11'b11110010110,
    11'b11101011101,
    11'b11101011100,
    11'b11101110000,
    11'b11110000011,
    11'b11101110010,
    11'b11101101010,
    11'b11110000110,
    11'b11110111000,
    11'b11110111101,
    11'b11110010011,
    11'b11101101010,
    11'b11101000001,
    11'b11100010110,
    11'b11011101011,
    11'b11011000000
};

parameter logic signed [`ACC_WIDTH-1:0] AZ_TEST_VECTOR[`NUM_ELEMENTS] = {
    11'b00011000100,
    11'b00011000110,
    11'b00011001010,
    11'b00011001111,
    11'b00011010100,
    11'b00011011001,
    11'b00011011101,
    11'b00011100101,
    11'b00011101100,
    11'b00011110100,
    11'b00011111010,
    11'b00011111011,
    11'b00011111101,
    11'b00011111110,
    11'b00011111110,
    11'b00011111110,
    11'b00011111101,
    11'b00100000000,
    11'b00100000011,
    11'b00100001010,
    11'b00100001111,
    11'b00100011010,
    11'b00100100100,
    11'b00100110011,
    11'b00101000001,
    11'b00101010100,
    11'b00101100100,
    11'b00101110100,
    11'b00110000010,
    11'b00110010010,
    11'b00110011010,
    11'b00110100010,
    11'b00110101000,
    11'b00110100110,
    11'b00110100100,
    11'b00110100011,
    11'b00110011001,
    11'b00110010110,
    11'b00110011100,
    11'b00110101000,
    11'b00110111100,
    11'b00111001001,
    11'b00111001101,
    11'b00111001001,
    11'b00110111001,
    11'b00110101100,
    11'b00110100001,
    11'b00110011010,
    11'b00110010011,
    11'b00110001111,
    11'b00110001101,
    11'b00110001011,
    11'b00110001010,
    11'b00110000110,
    11'b00110000101,
    11'b00110000101,
    11'b00110000110,
    11'b00110001010,
    11'b00110001101,
    11'b00110010110,
    11'b00110100000,
    11'b00110101100,
    11'b00110110110,
    11'b00111000100,
    11'b00111000100,
    11'b00110101111,
    11'b00110010110,
    11'b00101110110,
    11'b00101011101,
    11'b00101001010,
    11'b00101000111,
    11'b00101010110,
    11'b00101101111,
    11'b00110001110,
    11'b00110100111,
    11'b00110011101,
    11'b00101000011,
    11'b00100001110,
    11'b00010110010,
    11'b00001011000,
    11'b00000100100,
    11'b00010000000,
    11'b00100001001,
    11'b00111010101,
    11'b01010110011,
    11'b01101111000,
    11'b01110011110,
    11'b01101101110,
    11'b01011111010,
    11'b01000111011,
    11'b00110101100,
    11'b00100111000,
    11'b00011101101,
    11'b00011001000,
    11'b00011001111,
    11'b00011101101,
    11'b00100010001,
    11'b00100111000,
    11'b00101001000,
    11'b00101010000,
    11'b00101011100,
    11'b00101011100,
    11'b00101010011,
    11'b00101000100,
    11'b00101000100,
    11'b00101001011,
    11'b00101011010,
    11'b00101110001,
    11'b00110000000,
    11'b00110000110,
    11'b00110001110,
    11'b00110000011,
    11'b00101101111,
    11'b00101011011,
    11'b00101001100,
    11'b00101000011,
    11'b00101000110,
    11'b00101010000,
    11'b00101011111,
    11'b00101110111,
    11'b00110001010,
    11'b00110101100,
    11'b00111010110,
    11'b00111000001,
    11'b00110010000,
    11'b00110001011,
    11'b00110001111,
    11'b00110000101,
    11'b00101101010,
    11'b00101100010,
    11'b00101011000,
    11'b00101010001,
    11'b00101001000,
    11'b00101000111,
    11'b00101001011,
    11'b00101001000,
    11'b00101000001,
    11'b00100110000,
    11'b00100100011,
    11'b00100001000,
    11'b00011111000,
    11'b00011111010,
    11'b00100001001,
    11'b00100010011,
    11'b00100011101,
    11'b00100010011,
    11'b00100011100,
    11'b00100101010,
    11'b00100111100,
    11'b00101010001,
    11'b00101010101,
    11'b00101001000,
    11'b00101000011,
    11'b00100111111,
    11'b00100110100,
    11'b00100111011,
    11'b00100111010,
    11'b00101001010,
    11'b00101010010,
    11'b00101011001,
    11'b00101011010,
    11'b00101011010,
    11'b00101011100,
    11'b00101011111,
    11'b00101100011,
    11'b00101011101,
    11'b00101011111,
    11'b00101010111,
    11'b00101000110,
    11'b00101000010,
    11'b00101000101,
    11'b00101000100,
    11'b00101000000,
    11'b00101000011,
    11'b00101000111,
    11'b00101010011,
    11'b00110010110,
    11'b00110000001,
    11'b00101110001,
    11'b00101100111,
    11'b00101001011,
    11'b00100111111,
    11'b00100001111,
    11'b00100100001,
    11'b00100100011,
    11'b00011010100,
    11'b00001111010,
    11'b00000000100,
    11'b11101101000,
    11'b11101100001,
    11'b11110011101,
    11'b11111111101,
    11'b00001110111,
    11'b00011000110,
    11'b00100000010,
    11'b00100101011,
    11'b00101001001,
    11'b00101011100,
    11'b00101110110,
    11'b00110010100,
    11'b00111010011,
    11'b00111100111,
    11'b00110111011,
    11'b00110100110,
    11'b00110100011,
    11'b00101011011,
    11'b00100001101,
    11'b00011101111,
    11'b00010111010,
    11'b00010011010,
    11'b00010001101,
    11'b00010010011,
    11'b00010101000,
    11'b00011011000,
    11'b00100001010,
    11'b00101000101,
    11'b00110000001,
    11'b00111011000,
    11'b01000011110,
    11'b01001100001,
    11'b01010011100,
    11'b01011010111,
    11'b01011101111,
    11'b01011110100,
    11'b01011100100,
    11'b01010111110,
    11'b01001110100,
    11'b01000110101,
    11'b00111110111,
    11'b00110111110,
    11'b00101111111,
    11'b00101011100,
    11'b00100111111,
    11'b00100100111,
    11'b00100001101,
    11'b00011111100,
    11'b00011101111,
    11'b00011100010,
    11'b00011011100,
    11'b00011011001,
    11'b00011011000,
    11'b00011011010,
    11'b00011100001,
    11'b00011101101,
    11'b00011110011,
    11'b00010100100,
    11'b00001101111,
    11'b00100101110,
    11'b01001101111,
    11'b00101010000,
    11'b00010110111,
    11'b00011111100,
    11'b00101111100,
    11'b00100110100,
    11'b01000110011,
    11'b00110000011,
    11'b00100111010,
    11'b00100110110,
    11'b00101001101,
    11'b00100100011,
    11'b00100101101,
    11'b00100011111,
    11'b00100101000,
    11'b00100011110,
    11'b00100010111,
    11'b00100101100,
    11'b00100110110,
    11'b00100101100,
    11'b00100101100,
    11'b00100110011,
    11'b00100100011,
    11'b00100111011,
    11'b00100110110,
    11'b00100110100,
    11'b00100110110,
    11'b00100110101,
    11'b00100111110,
    11'b00100101001,
    11'b00100101101,
    11'b00100101111,
    11'b00100111001,
    11'b00100111111,
    11'b00100101111,
    11'b00100011000,
    11'b00100011111,
    11'b00100100010,
    11'b00100110111,
    11'b00100110100,
    11'b00100110100,
    11'b00100110100,
    11'b00100110011,
    11'b00100110000,
    11'b00100110000,
    11'b00100110011,
    11'b00100110001,
    11'b00100110001,
    11'b00100110001,
    11'b00100110001,
    11'b00100110001,
    11'b00100110001,
    11'b00100110000,
    11'b00100110001,
    11'b00100110000,
    11'b00100110000,
    11'b00100110000,
    11'b00100110000,
    11'b00100101111,
    11'b00100101111,
    11'b00100101111,
    11'b00100101111,
    11'b00100110000,
    11'b00100110000,
    11'b00100101111,
    11'b00100101111,
    11'b00100110001,
    11'b00100110001,
    11'b00100110010,
    11'b00100110010,
    11'b00100110011,
    11'b00100110011,
    11'b00100110010,
    11'b00100110001,
    11'b00100110010,
    11'b00100110001,
    11'b00100110001,
    11'b00100110001,
    11'b00100110001,
    11'b00100110001,
    11'b00100110001,
    11'b00100110001,
    11'b00100110001,
    11'b00100110001,
    11'b00100110001,
    11'b00100110001,
    11'b00100110010,
    11'b00100110010,
    11'b00100110000,
    11'b00100110001,
    11'b00100110001,
    11'b00100110010,
    11'b00100110011,
    11'b00100110100,
    11'b00100110100,
    11'b00100110010,
    11'b00100110011,
    11'b00100110100,
    11'b00100110011,
    11'b00100110001,
    11'b00100110001,
    11'b00100110001,
    11'b00100110010,
    11'b00100110011,
    11'b00100110011,
    11'b00100110100,
    11'b00100110011,
    11'b00100110001,
    11'b00100110001,
    11'b00100110010,
    11'b00100110010,
    11'b00100110010,
    11'b00100110010,
    11'b00100110001,
    11'b00100110001,
    11'b00100110010,
    11'b00100101111,
    11'b00100100000,
    11'b00100001011,
    11'b00100010100,
    11'b00100101100,
    11'b00100111100,
    11'b00101001000,
    11'b00101010010,
    11'b00101001000,
    11'b00100110011,
    11'b00101000100,
    11'b00100101100,
    11'b00100101101,
    11'b00100110001,
    11'b00100111010,
    11'b00100110110,
    11'b00100101110,
    11'b00100101010,
    11'b00100100110,
    11'b00100110010,
    11'b00100110110,
    11'b00100111010,
    11'b00100111100,
    11'b00100111000,
    11'b00100101110,
    11'b00100101111,
    11'b00100101111,
    11'b00100101111,
    11'b00100110111,
    11'b00100110100,
    11'b00100110000,
    11'b00100101100,
    11'b00100101100,
    11'b00100101111,
    11'b00100110100,
    11'b00100110110,
    11'b00100110111,
    11'b00100110111,
    11'b00100111000,
    11'b00100110110,
    11'b00100110110,
    11'b00101000110,
    11'b00110001000,
    11'b00111100111,
    11'b00110011111,
    11'b00100101100,
    11'b00100100110,
    11'b00011110111,
    11'b00101010010,
    11'b00111000101,
    11'b00110011010,
    11'b00101110001,
    11'b00101101111,
    11'b00100111000,
    11'b00101101010,
    11'b00101101000,
    11'b00100010101,
    11'b00010010110,
    11'b11101010011,
    11'b11110110110,
    11'b00001111010,
    11'b00001111001,
    11'b00000011100,
    11'b11111011101,
    11'b11110010000,
    11'b11110011011,
    11'b11111100110,
    11'b00100001110,
    11'b00110100001,
    11'b00100011111,
    11'b00011001001,
    11'b00001110000,
    11'b00100010111,
    11'b00100110011,
    11'b00101010100,
    11'b00101011101,
    11'b00101011111,
    11'b00110000001,
    11'b00101011101,
    11'b00101011111,
    11'b00101011100,
    11'b00101011001,
    11'b00101100001,
    11'b00101101100,
    11'b00101001111,
    11'b00100011000,
    11'b00011010011,
    11'b00010000011,
    11'b00001100110,
    11'b00001101101,
    11'b00010010010,
    11'b00011000111,
    11'b01001010101,
    11'b00110110011,
    11'b00110001111,
    11'b00110001101,
    11'b00101010101,
    11'b00101010110,
    11'b00101000110,
    11'b00101000010,
    11'b00101000100,
    11'b00101000100,
    11'b00101000011,
    11'b00101000110,
    11'b00101110010,
    11'b00110000011,
    11'b00101110100,
    11'b00101100011,
    11'b00100111010,
    11'b00100011000,
    11'b00011111111,
    11'b00011101100,
    11'b00011100011,
    11'b00011100110,
    11'b00011110000,
    11'b00011111101,
    11'b00110011101,
    11'b00101111100,
    11'b00101011011,
    11'b00101100001,
    11'b00101010011,
    11'b00101001101,
    11'b00101001010,
    11'b00101000110,
    11'b00101000001,
    11'b00101000001,
    11'b00101000000,
    11'b00100111111,
    11'b00101000110,
    11'b00101001100,
    11'b00101000011,
    11'b00101000000,
    11'b00100111011,
    11'b00100110001,
    11'b00100101011,
    11'b00100100100,
    11'b00100011011,
    11'b00100011001,
    11'b00100011100,
    11'b00101000111,
    11'b00101010101,
    11'b00101000100,
    11'b00101000110,
    11'b00100111011,
    11'b00100110110,
    11'b00100111101,
    11'b00100110011,
    11'b00100101001,
    11'b00100101111,
    11'b00100101000,
    11'b00100100011,
    11'b00101001110,
    11'b00101011001,
    11'b00101111011,
    11'b00101100011,
    11'b00111000110,
    11'b00011111101,
    11'b00101010011,
    11'b00100101110,
    11'b00011000011,
    11'b00001010010,
    11'b00001011010,
    11'b00111001010,
    11'b01001001111,
    11'b01011011100,
    11'b01001110101,
    11'b00110101001,
    11'b00101011111,
    11'b00110001010,
    11'b00111011010,
    11'b01000010010,
    11'b01000110001,
    11'b01001010101,
    11'b01001111001,
    11'b01001110000,
    11'b01000100110,
    11'b00110101000,
    11'b00100100000,
    11'b00011111000,
    11'b00011101000,
    11'b00011011100,
    11'b00011010110,
    11'b00011010101,
    11'b00011011100,
    11'b00011101100,
    11'b00100000110,
    11'b00100101100,
    11'b00101001010,
    11'b00101100110,
    11'b00110001110,
    11'b00110101101,
    11'b00111000100,
    11'b00111001000,
    11'b00111000011,
    11'b00110111100,
    11'b00110111010,
    11'b00110111110,
    11'b00111000011,
    11'b00110111110,
    11'b00110100001,
    11'b00101110101,
    11'b00101101100,
    11'b00110000111,
    11'b00110001100,
    11'b00110001111,
    11'b00110001110,
    11'b00110010011,
    11'b00110101001,
    11'b00110111110,
    11'b00111010110,
    11'b00111111011,
    11'b01000011001,
    11'b01000110100,
    11'b01000111110,
    11'b01000101111,
    11'b01000000111,
    11'b00111101000,
    11'b00111001111,
    11'b00111001111,
    11'b00111000111,
    11'b00111000001,
    11'b00110110110,
    11'b00110010100,
    11'b00101110010,
    11'b00101011100,
    11'b00101001100,
    11'b00100101011,
    11'b00001010100,
    11'b00000101110,
    11'b00001100010,
    11'b00100000011,
    11'b00101100011,
    11'b00110111000,
    11'b00111000011,
    11'b00110110100,
    11'b00111111010,
    11'b01001111100,
    11'b01010111100,
    11'b01010101010,
    11'b01011100001,
    11'b01010001100,
    11'b01000100010,
    11'b01000010010,
    11'b00100101101,
    11'b00110011001,
    11'b00111001100,
    11'b00110100101,
    11'b00101101100,
    11'b00100110001,
    11'b00011110101,
    11'b00010101100,
    11'b00001011011,
    11'b00000110001,
    11'b00000011000,
    11'b00000110110,
    11'b00001100001,
    11'b00000010110,
    11'b11110110011,
    11'b11101100011,
    11'b11100000001,
    11'b11010000110,
    11'b10111111001,
    11'b10110011100,
    11'b10110010001,
    11'b10110001101,
    11'b11100010110,
    11'b01110101011,
    11'b01111111111,
    11'b01111111111,
    11'b01111111111,
    11'b01111111111,
    11'b00101101101,
    11'b11011101111,
    11'b11010101100,
    11'b11101010011,
    11'b00001010110,
    11'b00101101101,
    11'b01001010101,
    11'b01001011011,
    11'b01000100001,
    11'b00110111010,
    11'b00011101100,
    11'b00000111110,
    11'b11110101010,
    11'b11101000110,
    11'b11100001101,
    11'b11011100110,
    11'b11011111111,
    11'b11101000111,
    11'b11110110110,
    11'b00001000100,
    11'b00010001111,
    11'b00010101111,
    11'b00011001001,
    11'b00011010001,
    11'b00010001000,
    11'b00001010000,
    11'b00000101000,
    11'b00000000100,
    11'b11110111000,
    11'b11101100100,
    11'b11100000110,
    11'b11011000001,
    11'b11010100100,
    11'b11010110110,
    11'b11011001000,
    11'b11011010100,
    11'b11011011001,
    11'b11011001110,
    11'b11011000111,
    11'b11011000001,
    11'b11010110011,
    11'b11010100011,
    11'b11010100010,
    11'b11010101000,
    11'b11010111100,
    11'b11011001101,
    11'b11011010010,
    11'b11011001000,
    11'b11011000110,
    11'b11011010001,
    11'b11011100011,
    11'b11011101001,
    11'b11011110100,
    11'b11011101010,
    11'b11011011010,
    11'b11011000111,
    11'b11010101001,
    11'b11010001100,
    11'b11001010100,
    11'b11000100100,
    11'b10111100010,
    11'b10110100001,
    11'b10101101111,
    11'b10101110001,
    11'b10110010110,
    11'b10111010010,
    11'b11000001101,
    11'b11001000010,
    11'b11001001100,
    11'b11000111100,
    11'b11000010110,
    11'b10111010011,
    11'b10110100100,
    11'b10110000110,
    11'b10101110100,
    11'b10101110000,
    11'b10101111011,
    11'b10110010001,
    11'b10110110010,
    11'b10111011010,
    11'b11000010101,
    11'b11001000010,
    11'b11001110111,
    11'b11010100110,
    11'b11011001100,
    11'b11011101100,
    11'b11100001000,
    11'b11100110100,
    11'b11101010100,
    11'b11101111010,
    11'b11110011101,
    11'b11111101010,
    11'b00000010011,
    11'b00000011000,
    11'b00000001001,
    11'b11111000101,
    11'b11100011010,
    11'b10101111100,
    11'b10111000010,
    11'b11000110010,
    11'b11001100110,
    11'b11010010001,
    11'b11010010001,
    11'b11010100001,
    11'b11011011011,
    11'b11110111010,
    11'b11110111101,
    11'b11101100000,
    11'b11100101001,
    11'b11100001011,
    11'b11100000010,
    11'b11100000110,
    11'b11100001010,
    11'b11100010001,
    11'b11100011000,
    11'b11100011000,
    11'b11100011100,
    11'b11100100000,
    11'b11100110100,
    11'b11101001010,
    11'b11101011000,
    11'b11101101001,
    11'b11110100011,
    11'b11110111101,
    11'b11111010000,
    11'b11111101001,
    11'b11111111010,
    11'b11111110001,
    11'b11111110011,
    11'b00000001111,
    11'b00000011100,
    11'b00000101101,
    11'b00000101010,
    11'b00001001000,
    11'b00001000101,
    11'b00001011001,
    11'b00001100110,
    11'b00001110011,
    11'b00010000100,
    11'b00010010111,
    11'b00010011000,
    11'b00010100100,
    11'b00010100011,
    11'b00010101011,
    11'b00010100011,
    11'b00010010001,
    11'b00001111011,
    11'b00010101011,
    11'b00010110011,
    11'b00011011000,
    11'b00011110011,
    11'b00100010001,
    11'b00100100011,
    11'b00011101111,
    11'b00010101111,
    11'b00010001111,
    11'b00001110001,
    11'b00001011011,
    11'b00001010101,
    11'b00001101010,
    11'b00010010100,
    11'b00011010000,
    11'b00011110011,
    11'b00100000101,
    11'b00100010001,
    11'b00100010110,
    11'b00100010110,
    11'b00100011010,
    11'b00100011100,
    11'b00100100011,
    11'b00100110100,
    11'b00101000001,
    11'b00101010111,
    11'b00101101000,
    11'b00101101010,
    11'b00101100011,
    11'b00101010010,
    11'b00101001100,
    11'b00101011000,
    11'b00100010111,
    11'b00101010001,
    11'b00101110110,
    11'b00101011100,
    11'b00101011001,
    11'b00101011111,
    11'b00100111100,
    11'b00101001010,
    11'b00100110011,
    11'b00100011101,
    11'b00100010011,
    11'b00100000011,
    11'b00011110001,
    11'b00011010011,
    11'b00010111011,
    11'b00010101000,
    11'b00010010010,
    11'b00010000001,
    11'b00001110001,
    11'b00001101010,
    11'b00001011011,
    11'b00001011010,
    11'b00001010011,
    11'b00001001111,
    11'b00001011000,
    11'b00001010100,
    11'b00001000101,
    11'b00000110100,
    11'b00000011100,
    11'b00000001111,
    11'b00000000001,
    11'b11111110101,
    11'b11111111000,
    11'b11111110101,
    11'b11111110001,
    11'b11111110101,
    11'b11111111010,
    11'b00000000001,
    11'b00000001010,
    11'b00000001100,
    11'b00000001111,
    11'b00000001101,
    11'b00000001101,
    11'b00000010110,
    11'b00000011000,
    11'b00000011010,
    11'b00000011010,
    11'b00000010000,
    11'b00000010010,
    11'b00000010000,
    11'b00000001000,
    11'b00000000000,
    11'b11111111100,
    11'b11111111010,
    11'b11111110011,
    11'b11111110111,
    11'b11111111100,
    11'b00000000000,
    11'b00000001000,
    11'b00000010100,
    11'b00000100101,
    11'b00000101101,
    11'b00000101001,
    11'b00000111100,
    11'b00001011010,
    11'b00000100111,
    11'b00000101000,
    11'b00010010000,
    11'b00010101111,
    11'b00010001101,
    11'b00010000000,
    11'b00011001111,
    11'b00011010101,
    11'b00011000101,
    11'b00011110101,
    11'b00010101010,
    11'b00100000001,
    11'b00101000101,
    11'b00100110110,
    11'b00100011110,
    11'b00100000010,
    11'b00001111001,
    11'b00100000100,
    11'b00011101010,
    11'b00001101111,
    11'b00010111000,
    11'b00010111000,
    11'b00011101110,
    11'b00011100001,
    11'b00100010001,
    11'b00101010110,
    11'b00101110100,
    11'b00111001101,
    11'b01000110011,
    11'b01000001101,
    11'b00110010110,
    11'b00101010010,
    11'b00101001111,
    11'b00001011010,
    11'b11101001111,
    11'b11101100000,
    11'b00001000110,
    11'b01000000101,
    11'b01111111111,
    11'b01111111111,
    11'b01111111111,
    11'b00111011111,
    11'b00110001000,
    11'b00100011111,
    11'b00000000011,
    11'b11101011101,
    11'b11100100110,
    11'b11111110001,
    11'b00011111010,
    11'b00111100110,
    11'b01001001101,
    11'b00111010001,
    11'b00110011111,
    11'b00110100001,
    11'b00111100100,
    11'b01011101111,
    11'b01001111010,
    11'b00111111011,
    11'b00111001010,
    11'b01001100100,
    11'b01101000000,
    11'b01111111111,
    11'b01111111111,
    11'b01111110011,
    11'b01110100001,
    11'b01101110110,
    11'b01100001111,
    11'b00111010100,
    11'b00101011011,
    11'b00111100011,
    11'b01010011101,
    11'b01100101010,
    11'b01101110000,
    11'b01111000101,
    11'b01111111111,
    11'b01111111111,
    11'b01111111111,
    11'b01100011111,
    11'b01001001011,
    11'b00010001010,
    11'b11110101000,
    11'b11101000100,
    11'b11101010001,
    11'b11111001100,
    11'b00001101011,
    11'b00011100011,
    11'b00100101101,
    11'b00101111111,
    11'b00110110101,
    11'b00111000011,
    11'b01000000100,
    11'b01001001101,
    11'b01000010010,
    11'b00111000110,
    11'b00100101011,
    11'b00011111100,
    11'b00001110011,
    11'b00001101100,
    11'b00000101111,
    11'b00000100111,
    11'b00000001101,
    11'b11111101001,
    11'b00001000000,
    11'b00010100110,
    11'b00011000111,
    11'b00010111101,
    11'b00010011101,
    11'b00010001000,
    11'b00010001000,
    11'b00001011000,
    11'b00000001000,
    11'b11110111101,
    11'b11111010011,
    11'b11111001000,
    11'b11110101000,
    11'b11111100011,
    11'b00000010110,
    11'b00000101000,
    11'b00000110100,
    11'b00001000010,
    11'b00001000110
};

parameter logic signed [`GYRO_WIDTH-1:0] WX_TEST_VECTOR[`NUM_ELEMENTS] = {
    14'b11111100011111,
    14'b11111100011100,
    14'b11111100010111,
    14'b11111100010010,
    14'b11111100001000,
    14'b11111011110110,
    14'b11111011100110,
    14'b11111011010010,
    14'b11111010111011,
    14'b11111010010111,
    14'b11111001111000,
    14'b11111001010111,
    14'b11111000110110,
    14'b11111000001010,
    14'b11110111101110,
    14'b11110111011010,
    14'b11110111001111,
    14'b11110111001101,
    14'b11110111010010,
    14'b11110111011111,
    14'b11110111110001,
    14'b11111000001111,
    14'b11111000100110,
    14'b11111000111011,
    14'b11111001001101,
    14'b11111001011111,
    14'b11111001100110,
    14'b11111001101100,
    14'b11111001101100,
    14'b11111001100100,
    14'b11111001011010,
    14'b11111001001101,
    14'b11111000110110,
    14'b11111000100110,
    14'b11111000010010,
    14'b11111000000101,
    14'b11111000001010,
    14'b11111000010111,
    14'b11111000101100,
    14'b11111001000000,
    14'b11111001001101,
    14'b11111001001101,
    14'b11111001001000,
    14'b11111001001000,
    14'b11111001001111,
    14'b11111001011111,
    14'b11111001110110,
    14'b11111010001101,
    14'b11111010110001,
    14'b11111011001101,
    14'b11111011101100,
    14'b11111100001010,
    14'b11111100110110,
    14'b11111101010111,
    14'b11111101111011,
    14'b11111110101001,
    14'b11111111001010,
    14'b11111111100100,
    14'b11111111110011,
    14'b00000000000000,
    14'b00000000000000,
    14'b11111111111101,
    14'b11111111111000,
    14'b11111111100110,
    14'b11111111001111,
    14'b11111110111101,
    14'b11111110111000,
    14'b11111111001010,
    14'b11111111101100,
    14'b00000000011111,
    14'b00000001011111,
    14'b00000010110011,
    14'b00000011011111,
    14'b00000011110001,
    14'b00000011101001,
    14'b00000010011111,
    14'b00000000110011,
    14'b11111110111011,
    14'b11111111001111,
    14'b00000000010100,
    14'b00000010111101,
    14'b00000111001010,
    14'b00001101010100,
    14'b00010001001000,
    14'b00010010101100,
    14'b00001111100110,
    14'b00001010001111,
    14'b00000100000011,
    14'b11111110110001,
    14'b11111010010111,
    14'b11111001011100,
    14'b11111010000011,
    14'b11111011100001,
    14'b11111101111011,
    14'b11111111100001,
    14'b00000000110011,
    14'b00000001110110,
    14'b00000010111011,
    14'b00000011100001,
    14'b00000011111101,
    14'b00000100100100,
    14'b00000101000101,
    14'b00000101100001,
    14'b00000101101110,
    14'b00000101101100,
    14'b00000101100100,
    14'b00000101001010,
    14'b00000100011111,
    14'b00000011101100,
    14'b00000010101100,
    14'b00000001101001,
    14'b00000000010100,
    14'b11111111101001,
    14'b11111111010100,
    14'b11111111010111,
    14'b11111111110001,
    14'b00000000001010,
    14'b00000000101001,
    14'b00000001000101,
    14'b00000001010111,
    14'b00000001010100,
    14'b00000000111000,
    14'b11111111001010,
    14'b11111110001111,
    14'b11111110000011,
    14'b11111101110011,
    14'b11111101011111,
    14'b11111101010010,
    14'b11111101001010,
    14'b11111100111101,
    14'b11111100111000,
    14'b11111100111101,
    14'b11111101010100,
    14'b11111101110001,
    14'b11111110000101,
    14'b11111110011100,
    14'b11111111000011,
    14'b11111111010111,
    14'b11111111011010,
    14'b11111111101110,
    14'b11111111110110,
    14'b11111111011100,
    14'b11111111000101,
    14'b11111111000011,
    14'b11111111000000,
    14'b11111111001101,
    14'b11111111010111,
    14'b11111110010111,
    14'b11111101001111,
    14'b11111100011111,
    14'b11111011111011,
    14'b11111011011111,
    14'b11111010111101,
    14'b11111010011111,
    14'b11111010001000,
    14'b11111010010010,
    14'b11111010000000,
    14'b11111001110011,
    14'b11111001100100,
    14'b11111001010111,
    14'b11111000111101,
    14'b11111000101100,
    14'b11111000010111,
    14'b11111000001101,
    14'b11111000001000,
    14'b11111000011010,
    14'b11111001000000,
    14'b11111001110011,
    14'b11111010100110,
    14'b11111011001010,
    14'b11111011101100,
    14'b11111100000101,
    14'b11111100010111,
    14'b11111100010111,
    14'b11111100001010,
    14'b11111011111011,
    14'b11111011100110,
    14'b11111011001010,
    14'b11111010101100,
    14'b11111010101100,
    14'b11111010110011,
    14'b11111010111000,
    14'b11111010001101,
    14'b11111001110110,
    14'b11111001010100,
    14'b11111001000101,
    14'b11111001100001,
    14'b11111010111000,
    14'b11111101101100,
    14'b11111110101001,
    14'b11111111101100,
    14'b00000000100100,
    14'b00000000100110,
    14'b11111111111011,
    14'b11111111001101,
    14'b11111110100110,
    14'b11111110001000,
    14'b11111101111000,
    14'b11111101101001,
    14'b11111101000000,
    14'b11111011101100,
    14'b11111011101110,
    14'b11111011110001,
    14'b11111010001000,
    14'b11111000010010,
    14'b11111000010111,
    14'b11110111110001,
    14'b11110111010010,
    14'b11111000100001,
    14'b11111001100001,
    14'b11111010010111,
    14'b11111011011010,
    14'b11111100100100,
    14'b11111110001101,
    14'b11111111110011,
    14'b00000001101110,
    14'b00000011101110,
    14'b00000101110001,
    14'b00000110101100,
    14'b00000110111101,
    14'b00000110100001,
    14'b00000100101100,
    14'b00000010101110,
    14'b00000000011111,
    14'b11111110010010,
    14'b11111100001101,
    14'b11111001111101,
    14'b11111000101110,
    14'b11110111111101,
    14'b11110111100001,
    14'b11110111010111,
    14'b11110111011111,
    14'b11110111101001,
    14'b11110111110110,
    14'b11111000001111,
    14'b11111000101001,
    14'b11111001001101,
    14'b11111010000101,
    14'b11111010110110,
    14'b11111011101100,
    14'b11111100100110,
    14'b11111101111011,
    14'b11111110111000,
    14'b11111111111000,
    14'b00000000100110,
    14'b11111110000101,
    14'b11111010111101,
    14'b11111010011100,
    14'b11111010100001,
    14'b11111001000011,
    14'b11110111110001,
    14'b11111000011010,
    14'b11110111000000,
    14'b11110110101100,
    14'b11110111111011,
    14'b11111010010100,
    14'b11111101001101,
    14'b11111110110001,
    14'b00000000000000,
    14'b00000000100001,
    14'b00000000110110,
    14'b00000000100110,
    14'b00000000001111,
    14'b00000000011010,
    14'b00000000010111,
    14'b00000000010010,
    14'b00000000001101,
    14'b00000000001101,
    14'b00000000001010,
    14'b00000000010010,
    14'b00000000001101,
    14'b11111111111101,
    14'b00000000000101,
    14'b00000000001010,
    14'b00000000001111,
    14'b00000000010100,
    14'b00000000010100,
    14'b00000000001010,
    14'b00000000001111,
    14'b00000000010010,
    14'b00000000001010,
    14'b11111111110011,
    14'b11111111011111,
    14'b11111111110110,
    14'b00000000010111,
    14'b00000000101100,
    14'b00000000111011,
    14'b00000000100100,
    14'b00000000011010,
    14'b00000000010111,
    14'b00000000010111,
    14'b00000000010111,
    14'b00000000011100,
    14'b00000000011010,
    14'b00000000010111,
    14'b00000000010111,
    14'b00000000010111,
    14'b00000000010100,
    14'b00000000010100,
    14'b00000000010100,
    14'b00000000010010,
    14'b00000000010010,
    14'b00000000010010,
    14'b00000000010010,
    14'b00000000010100,
    14'b00000000010100,
    14'b00000000010100,
    14'b00000000010100,
    14'b00000000010010,
    14'b00000000010010,
    14'b00000000010010,
    14'b00000000010010,
    14'b00000000010100,
    14'b00000000010111,
    14'b00000000010111,
    14'b00000000010111,
    14'b00000000010100,
    14'b00000000010100,
    14'b00000000010100,
    14'b00000000010100,
    14'b00000000010100,
    14'b00000000010100,
    14'b00000000010100,
    14'b00000000010100,
    14'b00000000010100,
    14'b00000000010100,
    14'b00000000010100,
    14'b00000000010100,
    14'b00000000010100,
    14'b00000000010100,
    14'b00000000010100,
    14'b00000000010100,
    14'b00000000010100,
    14'b00000000010100,
    14'b00000000010100,
    14'b00000000010100,
    14'b00000000010100,
    14'b00000000010100,
    14'b00000000010100,
    14'b00000000010100,
    14'b00000000010100,
    14'b00000000010100,
    14'b00000000010100,
    14'b00000000010100,
    14'b00000000010100,
    14'b00000000010100,
    14'b00000000010010,
    14'b00000000010010,
    14'b00000000010010,
    14'b00000000010010,
    14'b00000000010010,
    14'b00000000010010,
    14'b00000000010100,
    14'b00000000010100,
    14'b00000000010100,
    14'b00000000010100,
    14'b00000000010100,
    14'b00000000010100,
    14'b00000000010100,
    14'b00000000010100,
    14'b00000000010100,
    14'b00000000010100,
    14'b00000000010100,
    14'b00000000010100,
    14'b00000000010100,
    14'b00000000010010,
    14'b00000000001111,
    14'b00000000001101,
    14'b00000000001010,
    14'b00000000000101,
    14'b11111111111101,
    14'b11111111110011,
    14'b11111111111101,
    14'b00000000010100,
    14'b00000000110011,
    14'b00000000100110,
    14'b00000000011111,
    14'b00000000011111,
    14'b00000000011100,
    14'b00000000010111,
    14'b00000000010111,
    14'b00000000010010,
    14'b00000000010111,
    14'b00000000011010,
    14'b00000000011010,
    14'b00000000011010,
    14'b00000000010100,
    14'b00000000001101,
    14'b00000000001101,
    14'b00000000010010,
    14'b00000000010100,
    14'b00000000011010,
    14'b00000000011111,
    14'b00000000011100,
    14'b00000000011010,
    14'b00000000010111,
    14'b00000000010100,
    14'b00000000010100,
    14'b00000000010100,
    14'b00000000010100,
    14'b00000000010100,
    14'b00000000010100,
    14'b00000000010100,
    14'b00000000010100,
    14'b00000000010100,
    14'b00000000001111,
    14'b11111110101110,
    14'b11111011110011,
    14'b11111000000011,
    14'b11111000001101,
    14'b11111000101110,
    14'b11111010000101,
    14'b11111011011111,
    14'b11111101101100,
    14'b11111111100001,
    14'b00000001001101,
    14'b00000001110011,
    14'b00000001101110,
    14'b00000000000101,
    14'b11111111100001,
    14'b11111110001101,
    14'b11111011000011,
    14'b11110000110110,
    14'b11100110000011,
    14'b11101001110011,
    14'b11101101011010,
    14'b11110101011111,
    14'b11111111000000,
    14'b00001011000101,
    14'b00010100010111,
    14'b00011001001101,
    14'b00011011100100,
    14'b00010010111011,
    14'b00001010111011,
    14'b00000111100100,
    14'b00000111101100,
    14'b00000101110011,
    14'b00000100111011,
    14'b00000011010100,
    14'b00000010010010,
    14'b00000001010100,
    14'b00000000100110,
    14'b11111111100110,
    14'b11111110100100,
    14'b11111100011111,
    14'b11111011011010,
    14'b11111010000011,
    14'b11111000000000,
    14'b11110110110011,
    14'b11110110011100,
    14'b11110111100001,
    14'b11111011010010,
    14'b11111111011111,
    14'b00000100001000,
    14'b00001000011111,
    14'b00001011111011,
    14'b00001110000000,
    14'b00000111100001,
    14'b00000101000000,
    14'b00000100111000,
    14'b00000011000101,
    14'b00000000101001,
    14'b00000000101100,
    14'b00000000110011,
    14'b00000000101100,
    14'b00000000110001,
    14'b00000000100110,
    14'b00000000101001,
    14'b11111111110011,
    14'b11111110010100,
    14'b11111101001010,
    14'b11111100001111,
    14'b11111011101001,
    14'b11111011111011,
    14'b11111100101110,
    14'b11111101111101,
    14'b00000000000101,
    14'b00000001110011,
    14'b00000011011010,
    14'b00000100110011,
    14'b00000101111011,
    14'b00000011011100,
    14'b00000010111011,
    14'b00000010001010,
    14'b00000001011010,
    14'b00000001000011,
    14'b00000000110011,
    14'b00000000101001,
    14'b00000000100100,
    14'b00000000011100,
    14'b00000000011010,
    14'b00000000010111,
    14'b00000000001101,
    14'b11111111101001,
    14'b11111111011010,
    14'b11111111001111,
    14'b11111111001000,
    14'b11111111001010,
    14'b11111111010111,
    14'b11111111101100,
    14'b00000000010100,
    14'b00000000111101,
    14'b00000001100110,
    14'b00000010000101,
    14'b00000001010111,
    14'b00000001000101,
    14'b00000000110110,
    14'b00000000101100,
    14'b00000000100100,
    14'b00000000011100,
    14'b00000000011010,
    14'b00000000011111,
    14'b00000000100100,
    14'b00000000100110,
    14'b00000000101110,
    14'b00000000101001,
    14'b00000001000101,
    14'b00000001001010,
    14'b11111111000000,
    14'b11111100010111,
    14'b11111011010111,
    14'b11111101001000,
    14'b11111101010100,
    14'b11111110110110,
    14'b00000010111011,
    14'b00000110111101,
    14'b00001000111101,
    14'b00000111110110,
    14'b00001011101100,
    14'b00010001101001,
    14'b00010010101100,
    14'b00010001111101,
    14'b00010010001000,
    14'b00010101000101,
    14'b00010110001010,
    14'b00010010111000,
    14'b00001111001010,
    14'b00001100100001,
    14'b00001100110011,
    14'b00001110010111,
    14'b00010000110110,
    14'b00010100100110,
    14'b00010101111101,
    14'b00010101110110,
    14'b00010101001010,
    14'b00010011011100,
    14'b00010001111000,
    14'b00010000011111,
    14'b00001111011100,
    14'b00001110101110,
    14'b00001101110110,
    14'b00001101001000,
    14'b00001100010100,
    14'b00001011001010,
    14'b00001001110001,
    14'b00001001010100,
    14'b00001001000101,
    14'b00001000101110,
    14'b00001000010100,
    14'b00000111111011,
    14'b00000111010111,
    14'b00000110110110,
    14'b00000110100001,
    14'b00000110011111,
    14'b00000110001101,
    14'b00000101110001,
    14'b00000100110001,
    14'b00000100111000,
    14'b00000101100110,
    14'b00000101111000,
    14'b00000101101110,
    14'b00000101001111,
    14'b00000101001010,
    14'b00000100101100,
    14'b00000011011100,
    14'b00000010011100,
    14'b00000001011010,
    14'b00000000101001,
    14'b00000000101001,
    14'b00000001010100,
    14'b00000010001101,
    14'b00000011010010,
    14'b00000011111101,
    14'b00000100011111,
    14'b00000101000011,
    14'b00000101011111,
    14'b00000110001010,
    14'b00000110100001,
    14'b00000110010010,
    14'b00000110010111,
    14'b00000110011010,
    14'b00000010101110,
    14'b11111110010010,
    14'b11111110110011,
    14'b00000000010010,
    14'b00000001010100,
    14'b00000011001000,
    14'b00000100111011,
    14'b00000110001111,
    14'b00001000101001,
    14'b00001100010010,
    14'b00001110101110,
    14'b00001110000101,
    14'b00001110000011,
    14'b00001101001101,
    14'b00001001010111,
    14'b00001011001000,
    14'b00001010100110,
    14'b00001100000101,
    14'b00010000010010,
    14'b00010001110011,
    14'b00010001011111,
    14'b00001111110110,
    14'b00001111100001,
    14'b00001111011010,
    14'b00001111011111,
    14'b00001110011111,
    14'b00001110001101,
    14'b00001100111101,
    14'b00001011010111,
    14'b00001000100100,
    14'b00000110001101,
    14'b00000001100100,
    14'b11111011100001,
    14'b11110010000101,
    14'b11101100101110,
    14'b11101000111011,
    14'b11100111100100,
    14'b11101000111101,
    14'b11110010101100,
    14'b00001000000101,
    14'b00010001010111,
    14'b00001101000101,
    14'b00000110110110,
    14'b00000010111101,
    14'b00000100110001,
    14'b00001111101100,
    14'b00010111011111,
    14'b00011001000101,
    14'b00010101011010,
    14'b00001111110001,
    14'b00001001101001,
    14'b00001000111011,
    14'b00001000101110,
    14'b00001001111000,
    14'b00001110101001,
    14'b00010001101001,
    14'b00010010100001,
    14'b00010010101110,
    14'b00010011110110,
    14'b00010110000101,
    14'b00010111100100,
    14'b00011001000011,
    14'b00011010001111,
    14'b00011011100110,
    14'b00011100100100,
    14'b00011101101001,
    14'b00011110011111,
    14'b00011111000011,
    14'b00011101101001,
    14'b00011011101100,
    14'b00011010000101,
    14'b00011001001000,
    14'b00010111111101,
    14'b00010111001000,
    14'b00010110010111,
    14'b00010101110001,
    14'b00010101000011,
    14'b00010011110001,
    14'b00010010011100,
    14'b00010001000101,
    14'b00001111111011,
    14'b00001110001111,
    14'b00001101000000,
    14'b00001011101001,
    14'b00001010010100,
    14'b00001000101110,
    14'b00000111101100,
    14'b00000110101110,
    14'b00000110001000,
    14'b00000101110011,
    14'b00000101101001,
    14'b00000101100001,
    14'b00000101000101,
    14'b00000100111000,
    14'b00000100111101,
    14'b00000101010010,
    14'b00000101111101,
    14'b00000111000000,
    14'b00001001001101,
    14'b00001011001000,
    14'b00001101001101,
    14'b00001111010111,
    14'b00010001111011,
    14'b00010011011010,
    14'b00010100000101,
    14'b00010100000000,
    14'b00010011000101,
    14'b00010010000101,
    14'b00010001001010,
    14'b00010000010100,
    14'b00001111101001,
    14'b00001110111101,
    14'b00001110011100,
    14'b00001101101110,
    14'b00001100101100,
    14'b00001010110011,
    14'b00001001000011,
    14'b00000111000011,
    14'b00000100111101,
    14'b00000010111101,
    14'b00000000100001,
    14'b11111110111000,
    14'b11111101100100,
    14'b11111100011100,
    14'b11111010111000,
    14'b11111001010111,
    14'b11110111101001,
    14'b11110101101001,
    14'b11110010101110,
    14'b11110000110011,
    14'b11101110110011,
    14'b11101100110011,
    14'b11101011100110,
    14'b11101010110001,
    14'b11101010010111,
    14'b11101011110001,
    14'b11101101011111,
    14'b11101111011111,
    14'b11110001111101,
    14'b11110100100001,
    14'b11110110100110,
    14'b11101111001000,
    14'b11101100000000,
    14'b11101010001010,
    14'b11101001110011,
    14'b11101001110001,
    14'b11101001110110,
    14'b11101001011100,
    14'b11101001000101,
    14'b11101010111000,
    14'b11110000001010,
    14'b11110010101100,
    14'b11110011110110,
    14'b11110100001010,
    14'b11110011111011,
    14'b11110011110001,
    14'b11110011110011,
    14'b11110011100001,
    14'b11110011100100,
    14'b11110011101110,
    14'b11110011110011,
    14'b11110011011111,
    14'b11110011000011,
    14'b11110010000101,
    14'b11110000111000,
    14'b11101111110011,
    14'b11101110110001,
    14'b11101101100001,
    14'b11101100001111,
    14'b11101010111000,
    14'b11101001011010,
    14'b11100111100100,
    14'b11100101101100,
    14'b11100010110110,
    14'b11100000010111,
    14'b11011110010010,
    14'b11011101000101,
    14'b11011101000101,
    14'b11011101000101,
    14'b11011101000101,
    14'b11011101000101,
    14'b11011101000101,
    14'b11011101000101,
    14'b11011101000101,
    14'b11011101000101,
    14'b11011101000101,
    14'b11011101000101,
    14'b11011101000101,
    14'b11011101000101,
    14'b11011101000101,
    14'b11011110000000,
    14'b11100010001000,
    14'b11100101111101,
    14'b11101001011111,
    14'b11101100011111,
    14'b11101111011100,
    14'b11110010101100,
    14'b11110100010111,
    14'b11110100110011,
    14'b11110100011100,
    14'b11110011101100,
    14'b11110010001111,
    14'b11110000111101,
    14'b11101111101001,
    14'b11101110001111,
    14'b11101100011100,
    14'b11101011000000,
    14'b11101001011010,
    14'b11100111100100,
    14'b11100101011010,
    14'b11100010001000,
    14'b11011111010111,
    14'b11011101000101,
    14'b11011101000101,
    14'b11011101000101,
    14'b11011101000101,
    14'b11011101000101,
    14'b11011101000101,
    14'b11011101000101,
    14'b11011101000101,
    14'b11011101000101,
    14'b11011101000101,
    14'b11011101000101,
    14'b11011101000101,
    14'b11011101000101,
    14'b11011101000101,
    14'b11011101000101,
    14'b11011101000101,
    14'b11011101000101,
    14'b11011101000101,
    14'b11011101000101,
    14'b11011101000101,
    14'b11011101000101,
    14'b11011110110011,
    14'b11100001001000,
    14'b11100011010100,
    14'b11100101111101,
    14'b11100111110001,
    14'b11101001001000,
    14'b11101010001010,
    14'b11101011000011,
    14'b11101011011100,
    14'b11101011100100,
    14'b11101011100001,
    14'b11101011010111,
    14'b11101010111011,
    14'b11101010001101,
    14'b11101001001101,
    14'b11101000000101,
    14'b11100110100110,
    14'b11100101100110,
    14'b11100100110110,
    14'b11100100010100,
    14'b11100100001111,
    14'b11100100101110,
    14'b11100101011111,
    14'b11100110100100,
    14'b11100111110001,
    14'b11101001100100,
    14'b11101011001000,
    14'b11101100101110,
    14'b11101110011100,
    14'b11110000110011,
    14'b11110010101001,
    14'b11110100011111,
    14'b11110110001010,
    14'b11111000100001,
    14'b11111010001111,
    14'b11111011111011,
    14'b11111101100001,
    14'b11111111000000,
    14'b00000000111011,
    14'b00000010010010,
    14'b00000011101100,
    14'b00000101000101,
    14'b00000111000011,
    14'b00001000100100,
    14'b00001010000101,
    14'b00001011101110,
    14'b00001101011010,
    14'b00001111100100,
    14'b00010001000101,
    14'b00010010011111,
    14'b00010011110011,
    14'b00010101011010,
    14'b00010110100001,
    14'b00010111101110,
    14'b00011000101110,
    14'b00011001110110,
    14'b00011011001000,
    14'b00011011100001,
    14'b00011011011111,
    14'b00011011000011,
    14'b00011011010111,
    14'b00011011100001,
    14'b00011011000101,
    14'b00011010101110,
    14'b00011010010010,
    14'b00011001111000,
    14'b00011001111101,
    14'b00011000110110,
    14'b00011000000011,
    14'b00010111101110,
    14'b00011000000011,
    14'b00011001111000,
    14'b00011011011111,
    14'b00011011111101,
    14'b00011100110011,
    14'b00011110110110,
    14'b00100001100110,
    14'b00100010111011,
    14'b00100010111011,
    14'b00100010111011,
    14'b00100010111011,
    14'b00100010111011,
    14'b00100001111011,
    14'b00011111011010,
    14'b00011100000011,
    14'b00011010011010,
    14'b00011010010100,
    14'b00011011110110,
    14'b00100010111011,
    14'b00100010111011,
    14'b00100010111011,
    14'b00100010111011,
    14'b00100010111011,
    14'b00100010111011,
    14'b00100001100001,
    14'b00010111011010,
    14'b00010010001000,
    14'b00001110101110,
    14'b00001010100001,
    14'b00001011100110,
    14'b00001010010111,
    14'b00000110110011,
    14'b11111111001101,
    14'b11111110000101,
    14'b11111110100100,
    14'b00000001100001,
    14'b00000010111000,
    14'b11111111000101,
    14'b11110111011111,
    14'b11110000011010,
    14'b11101101110001,
    14'b11110100110001,
    14'b11110011111101,
    14'b11110010011010,
    14'b11110010101100,
    14'b11110100110110,
    14'b11110111011100,
    14'b11111010000101,
    14'b11111101001010,
    14'b11111111000101,
    14'b00000000110110,
    14'b00000001100110,
    14'b11111110100100,
    14'b11111010101100,
    14'b11110111001010,
    14'b11110100001010,
    14'b11110000101100,
    14'b11101101101110,
    14'b11101001110001,
    14'b11100101001111,
    14'b11011111000011,
    14'b11011101000101,
    14'b11011110011010,
    14'b11101101110011,
    14'b11111010001101,
    14'b11111011101001,
    14'b11111011011010,
    14'b11111101111000,
    14'b11111111100001,
    14'b11111111101001,
    14'b11111110000011,
    14'b11111101000011,
    14'b11111101111011,
    14'b11111100010111,
    14'b11111001000000,
    14'b11110011100100,
    14'b11101111110110,
    14'b11101101001000,
    14'b11101100100110,
    14'b11101011111000,
    14'b11101100011010,
    14'b11101110010111,
    14'b11110001010100,
    14'b11110100100110,
    14'b11110101110110,
    14'b11110100010100,
    14'b11101111111101,
    14'b11101101101110,
    14'b11110000111011,
    14'b11110011110110,
    14'b11110101110110,
    14'b11110111000101,
    14'b11110111110001,
    14'b11111000110001,
    14'b11111001111011,
    14'b11111010101001,
    14'b11111010011111,
    14'b11111010111101,
    14'b11111100011010,
    14'b11111101000000,
    14'b00000000000011,
    14'b00000000011111,
    14'b00000000101110,
    14'b00000000110011,
    14'b00000000110011,
    14'b00000000110001
};

parameter logic signed [`GYRO_WIDTH-1:0] WY_TEST_VECTOR[`NUM_ELEMENTS] = {
    14'b00000001011100,
    14'b00000001010010,
    14'b00000001001101,
    14'b00000001001000,
    14'b00000001000011,
    14'b00000000111101,
    14'b00000000111000,
    14'b00000000110110,
    14'b00000000110011,
    14'b00000000101110,
    14'b00000000101001,
    14'b00000000100100,
    14'b00000000011100,
    14'b00000000010010,
    14'b00000000001010,
    14'b00000000000011,
    14'b11111111111000,
    14'b11111111101110,
    14'b11111111100110,
    14'b11111111011111,
    14'b11111111010111,
    14'b11111111001111,
    14'b11111111001000,
    14'b11111111000011,
    14'b11111110111101,
    14'b11111110111011,
    14'b11111110111101,
    14'b11111111000000,
    14'b11111111000011,
    14'b11111111001000,
    14'b11111111001101,
    14'b11111111010010,
    14'b11111111010111,
    14'b11111111011100,
    14'b11111111100100,
    14'b11111111101001,
    14'b11111111101110,
    14'b11111111110110,
    14'b11111111111101,
    14'b11111111111101,
    14'b11111111111011,
    14'b11111111110110,
    14'b11111111101100,
    14'b11111111100001,
    14'b11111111010111,
    14'b11111111001111,
    14'b11111111001010,
    14'b11111111001000,
    14'b11111111001000,
    14'b11111111001010,
    14'b11111111001111,
    14'b11111111010100,
    14'b11111111011100,
    14'b11111111100001,
    14'b11111111100110,
    14'b11111111101110,
    14'b11111111110110,
    14'b11111111111011,
    14'b11111111111101,
    14'b00000000000011,
    14'b00000000000101,
    14'b00000000001010,
    14'b00000000001101,
    14'b00000000001101,
    14'b00000000000011,
    14'b11111111110011,
    14'b11111111101110,
    14'b11111111100110,
    14'b11111111100001,
    14'b11111111100100,
    14'b11111111101110,
    14'b11111111111000,
    14'b00000000000011,
    14'b00000000001000,
    14'b00000000001010,
    14'b00000000010111,
    14'b00000000111101,
    14'b00000001111000,
    14'b00000010110110,
    14'b00000100001111,
    14'b00000110011111,
    14'b00000111101100,
    14'b00001000001000,
    14'b00001000000101,
    14'b00000110111011,
    14'b00000100111000,
    14'b00000011001010,
    14'b00000001011111,
    14'b00000000000011,
    14'b11111110110001,
    14'b11111110010100,
    14'b11111110011100,
    14'b11111111000000,
    14'b11111111111101,
    14'b00000000101110,
    14'b00000001010111,
    14'b00000001111011,
    14'b00000010010111,
    14'b00000010100100,
    14'b00000010101001,
    14'b00000010100100,
    14'b00000010010100,
    14'b00000001111000,
    14'b00000001101100,
    14'b00000001100001,
    14'b00000001010100,
    14'b00000001000011,
    14'b00000000111011,
    14'b00000000101001,
    14'b00000000011111,
    14'b00000000010111,
    14'b00000000001101,
    14'b00000000001010,
    14'b00000000010010,
    14'b00000000011010,
    14'b00000000100100,
    14'b00000000100110,
    14'b00000000101001,
    14'b00000000100110,
    14'b00000000011111,
    14'b00000000010100,
    14'b00000000001101,
    14'b00000000000011,
    14'b11111111101100,
    14'b11111111100100,
    14'b11111111101100,
    14'b11111111110001,
    14'b11111111110001,
    14'b11111111101100,
    14'b11111111101001,
    14'b11111111100100,
    14'b11111111100001,
    14'b11111111011010,
    14'b11111111010100,
    14'b11111111001010,
    14'b11111111000011,
    14'b11111110110110,
    14'b11111110110110,
    14'b11111111000000,
    14'b11111111001010,
    14'b11111111100100,
    14'b00000000000000,
    14'b00000000010111,
    14'b00000000100100,
    14'b00000000110001,
    14'b00000000110110,
    14'b00000000111101,
    14'b00000001000101,
    14'b00000001001000,
    14'b00000000110001,
    14'b00000000001101,
    14'b11111111101001,
    14'b11111111010010,
    14'b11111110100110,
    14'b11111110100001,
    14'b11111110010100,
    14'b11111110011010,
    14'b11111110100001,
    14'b11111110100110,
    14'b11111110101100,
    14'b11111110101110,
    14'b11111110110011,
    14'b11111110111101,
    14'b11111111010010,
    14'b11111111011111,
    14'b11111111100100,
    14'b11111111101001,
    14'b11111111100001,
    14'b11111111011100,
    14'b11111111100001,
    14'b11111111101100,
    14'b11111111110011,
    14'b00000000000000,
    14'b00000000001000,
    14'b00000000001010,
    14'b00000000001101,
    14'b11111110010111,
    14'b11111101000000,
    14'b11111100010010,
    14'b11111011110011,
    14'b11111011110110,
    14'b11111011110011,
    14'b11111011111000,
    14'b11111100100001,
    14'b11111011100001,
    14'b11111011001010,
    14'b11111011100001,
    14'b11111100001000,
    14'b11111110100001,
    14'b00000001000000,
    14'b00000011001101,
    14'b00000100110110,
    14'b00000110010100,
    14'b00000111000011,
    14'b00000111011100,
    14'b00000111101100,
    14'b00000111101100,
    14'b00000111101110,
    14'b00000111100100,
    14'b00000111011111,
    14'b00000111000000,
    14'b00000101111011,
    14'b00000101000000,
    14'b00000100101110,
    14'b00000100001000,
    14'b00000011101100,
    14'b00000100001101,
    14'b00000101001101,
    14'b00000110011010,
    14'b00000111100001,
    14'b00001000101110,
    14'b00001001110011,
    14'b00001010110011,
    14'b00001100001000,
    14'b00001101000000,
    14'b00001101100100,
    14'b00001101111000,
    14'b00001101111011,
    14'b00001101101001,
    14'b00001101000101,
    14'b00001100010010,
    14'b00001010110011,
    14'b00001001010111,
    14'b00000111101100,
    14'b00000101110011,
    14'b00000011111011,
    14'b00000001100001,
    14'b11111111111000,
    14'b11111110011100,
    14'b11111101001010,
    14'b11111011110001,
    14'b11111010111011,
    14'b11111010010100,
    14'b11111001111101,
    14'b11111001110011,
    14'b11111001111011,
    14'b11111010010010,
    14'b11111011000101,
    14'b11111011111000,
    14'b11111100110001,
    14'b11111101110001,
    14'b11111111000101,
    14'b00000000000101,
    14'b00000001000011,
    14'b00000001110011,
    14'b00000010000101,
    14'b00000010011010,
    14'b00000010100110,
    14'b00000001011100,
    14'b11111111001010,
    14'b11111111101100,
    14'b11111111011111,
    14'b11111110101110,
    14'b11111100111101,
    14'b11111010100001,
    14'b11111001110001,
    14'b11111001100100,
    14'b11111010001101,
    14'b11111011010010,
    14'b11111011101110,
    14'b11111011101001,
    14'b11111011111101,
    14'b11111100110001,
    14'b11111101101100,
    14'b11111110111011,
    14'b00000000000101,
    14'b00000000111101,
    14'b00000000111101,
    14'b00000000110110,
    14'b00000000011010,
    14'b00000000001111,
    14'b00000000001101,
    14'b11111111111000,
    14'b11111111100100,
    14'b11111111000101,
    14'b11111110010111,
    14'b11111101111101,
    14'b11111101110011,
    14'b11111101101110,
    14'b11111101111000,
    14'b11111110000011,
    14'b11111110001111,
    14'b11111110011111,
    14'b11111111000000,
    14'b11111111011100,
    14'b11111111111000,
    14'b00000000010111,
    14'b00000000110001,
    14'b00000000111000,
    14'b00000000111101,
    14'b00000000111101,
    14'b00000000111011,
    14'b00000000110011,
    14'b00000000101001,
    14'b00000000011010,
    14'b00000000000101,
    14'b11111111100110,
    14'b11111111010100,
    14'b11111111000101,
    14'b11111110111011,
    14'b11111110110011,
    14'b11111110110001,
    14'b11111110101110,
    14'b11111110110001,
    14'b11111110111011,
    14'b11111111000101,
    14'b11111111010100,
    14'b11111111100001,
    14'b11111111110011,
    14'b11111111111101,
    14'b00000000001000,
    14'b00000000001101,
    14'b00000000010100,
    14'b00000000010111,
    14'b00000000010111,
    14'b00000000010010,
    14'b00000000001010,
    14'b00000000000000,
    14'b11111111110110,
    14'b11111111101110,
    14'b11111111100110,
    14'b11111111011100,
    14'b11111111010100,
    14'b11111111010010,
    14'b11111111001111,
    14'b11111111001111,
    14'b11111111010010,
    14'b11111111010100,
    14'b11111111011100,
    14'b11111111100100,
    14'b11111111101001,
    14'b11111111110001,
    14'b11111111111000,
    14'b11111111111101,
    14'b00000000000000,
    14'b00000000000011,
    14'b00000000000011,
    14'b00000000000000,
    14'b11111111111101,
    14'b11111111111011,
    14'b11111111110110,
    14'b11111111110001,
    14'b11111111101100,
    14'b11111111101001,
    14'b11111111100100,
    14'b11111111100001,
    14'b11111111100001,
    14'b11111111011111,
    14'b11111111100001,
    14'b11111111100001,
    14'b11111111100100,
    14'b11111111100110,
    14'b11111111101100,
    14'b11111111101110,
    14'b11111111110001,
    14'b11111111110110,
    14'b11111111111000,
    14'b11111111111000,
    14'b11111111111000,
    14'b11111111111000,
    14'b11111111111000,
    14'b11111111110110,
    14'b11111111110011,
    14'b11111111110011,
    14'b11111111101110,
    14'b11111111101110,
    14'b11111111101110,
    14'b11111111110001,
    14'b11111111111000,
    14'b11111111110110,
    14'b11111111110011,
    14'b00000000001000,
    14'b00000000010100,
    14'b00000000100001,
    14'b00000000111011,
    14'b00000001001000,
    14'b00000000111011,
    14'b00000000010111,
    14'b11111111100100,
    14'b11111110111101,
    14'b11111110101100,
    14'b11111110101100,
    14'b11111110101110,
    14'b11111110101110,
    14'b11111110100001,
    14'b11111110011010,
    14'b11111110011010,
    14'b11111110100110,
    14'b11111111000101,
    14'b11111111011010,
    14'b11111111101100,
    14'b11111111110110,
    14'b11111111111011,
    14'b00000000000000,
    14'b00000000001000,
    14'b00000000001111,
    14'b00000000010111,
    14'b00000000010111,
    14'b00000000010010,
    14'b00000000001000,
    14'b11111111111000,
    14'b11111111101110,
    14'b11111111100110,
    14'b11111111100001,
    14'b11111111011100,
    14'b11111111001010,
    14'b11111111101001,
    14'b11111111101001,
    14'b11111110111000,
    14'b11111101011100,
    14'b11111100110001,
    14'b11111011010111,
    14'b11111100100110,
    14'b11111100011111,
    14'b11111011101001,
    14'b11111010100110,
    14'b11111001100100,
    14'b11111000111000,
    14'b11111001001111,
    14'b11111001110110,
    14'b11111010110001,
    14'b11111100010100,
    14'b11111111101001,
    14'b00000010000101,
    14'b11111101011111,
    14'b11111101010100,
    14'b11111110011100,
    14'b00000001001010,
    14'b00000100010100,
    14'b00001000111000,
    14'b00001100000011,
    14'b00001100100100,
    14'b00001000111011,
    14'b00000111101110,
    14'b00000101001111,
    14'b00000010110011,
    14'b00000001010100,
    14'b00000001100100,
    14'b11111111101001,
    14'b11111100110110,
    14'b11111001100110,
    14'b11110111001000,
    14'b11110101011100,
    14'b11110101011111,
    14'b11110110100100,
    14'b11110111010111,
    14'b11111000100100,
    14'b11111010001000,
    14'b11111011100001,
    14'b11111101010100,
    14'b11111111100001,
    14'b00000010101001,
    14'b00000100111011,
    14'b00000110111101,
    14'b00001000011111,
    14'b00001001011111,
    14'b00001000101100,
    14'b00001001010010,
    14'b00001000000101,
    14'b00000110010111,
    14'b00000100010010,
    14'b00000011101001,
    14'b00000001110011,
    14'b11111111111101,
    14'b11111110000000,
    14'b11111100100100,
    14'b11111011001111,
    14'b11111010100001,
    14'b11111010000000,
    14'b11111001110011,
    14'b11111001111011,
    14'b11111010001101,
    14'b11111010111000,
    14'b11111011111000,
    14'b11111101001000,
    14'b11111110011100,
    14'b00000000001000,
    14'b00000001010010,
    14'b00000010001111,
    14'b00000011000011,
    14'b00000011101100,
    14'b00000011110001,
    14'b00000011111011,
    14'b00000011010100,
    14'b00000010100001,
    14'b00000010000101,
    14'b00000001011010,
    14'b00000000101001,
    14'b00000000000011,
    14'b11111111001000,
    14'b11111110011010,
    14'b11111101111011,
    14'b11111101101001,
    14'b11111101011010,
    14'b11111101011100,
    14'b11111101101001,
    14'b11111101110110,
    14'b11111110010111,
    14'b11111110110110,
    14'b11111111010111,
    14'b00000000001000,
    14'b00000000101001,
    14'b00000001001000,
    14'b00000001011010,
    14'b00000001100001,
    14'b00000001100110,
    14'b00000001011010,
    14'b00000001001010,
    14'b00000001000000,
    14'b00000000101100,
    14'b00000000011010,
    14'b00000000000011,
    14'b11111111101100,
    14'b11111111011100,
    14'b11111111001010,
    14'b11111110000101,
    14'b11111000000011,
    14'b11110001000101,
    14'b11111001001010,
    14'b11111011011010,
    14'b11111100101001,
    14'b11111100100001,
    14'b11111101100100,
    14'b11111111001111,
    14'b00000100000011,
    14'b00001000001010,
    14'b00001010011010,
    14'b00001010011111,
    14'b00001001101110,
    14'b00000111001101,
    14'b00000111010100,
    14'b00001001010100,
    14'b00001010100100,
    14'b00001010010100,
    14'b00001001011010,
    14'b00000111100110,
    14'b00000101110110,
    14'b00000011100001,
    14'b00000001101110,
    14'b11111111101110,
    14'b11111101110011,
    14'b11111100101001,
    14'b11111100011111,
    14'b11111100101100,
    14'b11111101010100,
    14'b11111110011100,
    14'b11111111001111,
    14'b00000000000000,
    14'b00000000101001,
    14'b00000001001101,
    14'b00000001111000,
    14'b00000010001111,
    14'b00000010011100,
    14'b00000010011010,
    14'b00000001100110,
    14'b00000000110110,
    14'b00000000000011,
    14'b11111111010010,
    14'b11111110011100,
    14'b11111101011111,
    14'b11111100110001,
    14'b11111100000101,
    14'b11111011010111,
    14'b11111010101110,
    14'b11111010010100,
    14'b11111010010100,
    14'b11111010011010,
    14'b11111010001000,
    14'b11111001111000,
    14'b11111001101110,
    14'b11111001101100,
    14'b11111001101001,
    14'b11111001011010,
    14'b11111001001111,
    14'b11111001000000,
    14'b11111000011111,
    14'b11110111110011,
    14'b11110110100110,
    14'b11110101101001,
    14'b11110100110001,
    14'b11110100001000,
    14'b11110011011010,
    14'b11110010111011,
    14'b11110010010111,
    14'b11110001111101,
    14'b11110001011111,
    14'b11110000111000,
    14'b11110000101100,
    14'b11110000101110,
    14'b11110000111000,
    14'b11110001001101,
    14'b11110010110110,
    14'b11110101001111,
    14'b11110111010111,
    14'b11111000011010,
    14'b11111000101001,
    14'b11110111111000,
    14'b11110110111000,
    14'b11110110000000,
    14'b11110101010100,
    14'b11110100000011,
    14'b11110010000101,
    14'b11110000101001,
    14'b11101110011100,
    14'b11101100011111,
    14'b11101011110001,
    14'b11101011000000,
    14'b11101010100110,
    14'b11101010101110,
    14'b11101001111000,
    14'b11101001011100,
    14'b11101001101110,
    14'b11101001111000,
    14'b11101010010010,
    14'b11101010011010,
    14'b11101011010100,
    14'b11101100101110,
    14'b11101101101100,
    14'b11101110110001,
    14'b11101111000011,
    14'b11101101100100,
    14'b11101100110110,
    14'b11101011111000,
    14'b11101010011111,
    14'b11100111001111,
    14'b11100100101110,
    14'b11100100001111,
    14'b11100100011100,
    14'b11100101111011,
    14'b11101110101100,
    14'b11111010000011,
    14'b11111000111011,
    14'b11110110110110,
    14'b11110011001111,
    14'b11101110111011,
    14'b11101110010100,
    14'b11110011010100,
    14'b11110111011010,
    14'b11111001111000,
    14'b11111010100100,
    14'b11111001110011,
    14'b11110111000011,
    14'b11110100011100,
    14'b11110010001111,
    14'b11110000001111,
    14'b11101110001111,
    14'b11101110000011,
    14'b11101111001010,
    14'b11110001001010,
    14'b11110011100001,
    14'b11110110111101,
    14'b11111001101100,
    14'b11111100000000,
    14'b11111101100100,
    14'b11111110001101,
    14'b11111101110001,
    14'b11111100111000,
    14'b11111011111000,
    14'b11111001111101,
    14'b11110111011111,
    14'b11110110001111,
    14'b11110101011111,
    14'b11110100111011,
    14'b11110100001111,
    14'b11110011111011,
    14'b11110100001010,
    14'b11110100110001,
    14'b11110101100001,
    14'b11110110011100,
    14'b11110110111011,
    14'b11110111011010,
    14'b11110111101110,
    14'b11110111111101,
    14'b11111000000000,
    14'b11110111111011,
    14'b11110111110011,
    14'b11110111101110,
    14'b11110111101001,
    14'b11110111011111,
    14'b11110111001111,
    14'b11110110111000,
    14'b11110110011100,
    14'b11110110001101,
    14'b11110110010010,
    14'b11110110011111,
    14'b11110111000000,
    14'b11110111100110,
    14'b11111000010100,
    14'b11111000111000,
    14'b11111001111011,
    14'b11111010101001,
    14'b11111011011010,
    14'b11111100001010,
    14'b11111101010010,
    14'b11111110000101,
    14'b11111110111101,
    14'b11111111111101,
    14'b00000001011010,
    14'b00000010011100,
    14'b00000011001101,
    14'b00000011100100,
    14'b00000011011010,
    14'b00000010100001,
    14'b00000001100001,
    14'b00000000011100,
    14'b11111111011111,
    14'b11111110100001,
    14'b11111110001010,
    14'b11111110000011,
    14'b11111110001000,
    14'b11111110010100,
    14'b11111110101100,
    14'b11111111000000,
    14'b11111111010100,
    14'b11111111100100,
    14'b11111111101110,
    14'b11111111101001,
    14'b11111111011010,
    14'b11111111001010,
    14'b11111110110011,
    14'b11111110100100,
    14'b11111110010100,
    14'b11111110000000,
    14'b11111101100110,
    14'b11111101010010,
    14'b11111100100100,
    14'b11111010101110,
    14'b11111000111101,
    14'b11110110111000,
    14'b11110100011100,
    14'b11110001110110,
    14'b11110000000000,
    14'b11110101000000,
    14'b11110111010100,
    14'b11111001100110,
    14'b11111010100100,
    14'b11111011001010,
    14'b11111011001000,
    14'b11111010101100,
    14'b11111010001101,
    14'b11111001000011,
    14'b11110110000000,
    14'b11110100011010,
    14'b11110011100001,
    14'b11110011001010,
    14'b11110011001101,
    14'b11110011011100,
    14'b11110011111000,
    14'b11110100100100,
    14'b11110101001000,
    14'b11110101010111,
    14'b11110101011111,
    14'b11110101100110,
    14'b11110101101001,
    14'b11110101110001,
    14'b11110101111011,
    14'b11110110001000,
    14'b11110110001000,
    14'b11110110000011,
    14'b11110101111101,
    14'b11110101101100,
    14'b11110101011100,
    14'b11110101001101,
    14'b11110101000000,
    14'b11110100101110,
    14'b11110100011111,
    14'b11110100001101,
    14'b11110100001010,
    14'b11110100011100,
    14'b11110101001111,
    14'b11110110000101,
    14'b11110111000101,
    14'b11110111111101,
    14'b11111001000101,
    14'b11111001110110,
    14'b11111010101001,
    14'b11111011111000,
    14'b11111100111000,
    14'b11111111001101,
    14'b00000000101100,
    14'b00000001110001,
    14'b00000011001000,
    14'b00000100100100,
    14'b00000100101001,
    14'b00000100101110,
    14'b00000101010111,
    14'b00000110010111,
    14'b00001000001101,
    14'b00001001000000,
    14'b00001000111000,
    14'b00000111111000,
    14'b00000101111101,
    14'b00000010111011,
    14'b00000000101100,
    14'b11111111000011,
    14'b11111110001010,
    14'b11111110001111,
    14'b11111110101100,
    14'b11111111001010,
    14'b11111111100100,
    14'b11111111110011,
    14'b11111111110011,
    14'b11111111101100,
    14'b11111111100100,
    14'b11111111101100,
    14'b00000000001111,
    14'b00000000110110,
    14'b00000001011111,
    14'b00000010000101,
    14'b00000010110001,
    14'b00000011001010,
    14'b00000011101001,
    14'b00000100001010,
    14'b00000100011111,
    14'b00000101100100,
    14'b00000110011111,
    14'b00000110011010,
    14'b00000110001000,
    14'b00000110101110,
    14'b00000110001101,
    14'b00000110000101,
    14'b00000110100100,
    14'b00000110010010,
    14'b00000110000011,
    14'b00000101101100,
    14'b00000101001000,
    14'b00000100011100,
    14'b00000011101100,
    14'b00000011001010,
    14'b00000010110110,
    14'b00000010100110,
    14'b00000010011111,
    14'b00000010010111,
    14'b00000010001111,
    14'b00000010001010,
    14'b00000010001000,
    14'b00000001111011,
    14'b00000001111011,
    14'b00000010000101,
    14'b00000010001010,
    14'b00000010011010,
    14'b00000010101001,
    14'b00000010110110,
    14'b00000011001010,
    14'b00000011010010,
    14'b00000011011010,
    14'b00000011010111,
    14'b00000011001000,
    14'b00000010111011,
    14'b00000010101001,
    14'b00000010010100,
    14'b00000010001000,
    14'b00000001111011,
    14'b00000001101110,
    14'b00000001101100,
    14'b00000001100100,
    14'b00000001100110,
    14'b00000001100110,
    14'b00000001011111,
    14'b00000001011010,
    14'b00000001010010,
    14'b00000001001101,
    14'b00000001001101,
    14'b00000001000101,
    14'b00000001000000,
    14'b00000000111011,
    14'b00000000110011,
    14'b00000000100110,
    14'b00000000011010,
    14'b00000000001010,
    14'b11111111110011,
    14'b11111111010100,
    14'b11111110111101,
    14'b11111110100110,
    14'b11111110010100,
    14'b11111110000011,
    14'b11111110001000,
    14'b11111110011111,
    14'b11111110101100,
    14'b11111111001010,
    14'b00000000101001,
    14'b00000000111101,
    14'b00000000101110,
    14'b00000000110011,
    14'b00000001010010,
    14'b00000001011010,
    14'b00000000111101,
    14'b00000001100001,
    14'b00000001100100,
    14'b00000001101001,
    14'b00000010100001,
    14'b00000001010111,
    14'b00000000101100,
    14'b00000000010010,
    14'b11111111111011,
    14'b00000001000000,
    14'b00000010001010,
    14'b00000010001101,
    14'b00000011011100,
    14'b00000101111000,
    14'b00001000000011,
    14'b00001001001010,
    14'b00001010111101,
    14'b00001100101100,
    14'b00001100011111,
    14'b00001011110001,
    14'b00001010110110,
    14'b00001000110011,
    14'b00000101110110,
    14'b00000100101100,
    14'b00000100011100,
    14'b00000100010111,
    14'b00000010101001,
    14'b00000010001000,
    14'b00000011110110,
    14'b00000101001111,
    14'b00000100100100,
    14'b00000111000101,
    14'b11111001001101,
    14'b11101111001000,
    14'b11101110010111,
    14'b11101110001000,
    14'b11101111110001,
    14'b11110001111000,
    14'b11110110011111,
    14'b11111011101110,
    14'b00000010000011,
    14'b00000100100001,
    14'b00000101001010,
    14'b00000100011100,
    14'b00000011010111,
    14'b00000011010100,
    14'b00000011101001,
    14'b00000011011010,
    14'b00000010100110,
    14'b11110111111000,
    14'b11110111101001,
    14'b11111000010100,
    14'b11111010011100,
    14'b11111011111000,
    14'b11111010110110,
    14'b11110111001101,
    14'b11110010011100,
    14'b11110000000101,
    14'b11101101101100,
    14'b11101011010111,
    14'b11101001100001,
    14'b11101010001101,
    14'b11101010111101,
    14'b11101010000101,
    14'b11100111011111,
    14'b11100101100001,
    14'b11100011100001,
    14'b11100001011010,
    14'b11011101001010,
    14'b11011101000101,
    14'b11011101000101,
    14'b11011101000101,
    14'b11011101000101,
    14'b11011101000101,
    14'b11011110000101,
    14'b11100100101110,
    14'b11101000010111,
    14'b11101010010100,
    14'b11101011001101,
    14'b11101011001010,
    14'b11101010101100,
    14'b11101001100110,
    14'b11101000011111,
    14'b11100110110001,
    14'b11100101011100,
    14'b11100011101001,
    14'b11100010100110,
    14'b11100010000101,
    14'b11100010110011,
    14'b11100010111101,
    14'b11100100000011,
    14'b11100100100110,
    14'b11100101100110,
    14'b11100110011010,
    14'b11100111101001,
    14'b11101001011010,
    14'b11101001011010,
    14'b11101000111000,
    14'b11101000100110,
    14'b11101000111101,
    14'b11101001100100,
    14'b11101010000101,
    14'b11101010110110,
    14'b11101011011100,
    14'b11101100111101,
    14'b11101110100110,
    14'b11101111100100,
    14'b11110001000011,
    14'b11110101100100,
    14'b11110110001101,
    14'b11110110010010,
    14'b11110110001111,
    14'b11110110000000,
    14'b11110101101100
};

parameter logic signed [`GYRO_WIDTH-1:0] WZ_TEST_VECTOR[`NUM_ELEMENTS] = {
    14'b11111101010100,
    14'b11111101001000,
    14'b11111101000011,
    14'b11111101000000,
    14'b11111100111011,
    14'b11111100110011,
    14'b11111100101001,
    14'b11111100011100,
    14'b11111100001101,
    14'b11111011110110,
    14'b11111011100100,
    14'b11111011001111,
    14'b11111010111011,
    14'b11111010100001,
    14'b11111010010010,
    14'b11111010000101,
    14'b11111001111011,
    14'b11111001110011,
    14'b11111001110110,
    14'b11111001111011,
    14'b11111010000101,
    14'b11111010010111,
    14'b11111010100100,
    14'b11111010110001,
    14'b11111010111101,
    14'b11111011001101,
    14'b11111011010111,
    14'b11111011011111,
    14'b11111011100110,
    14'b11111011110001,
    14'b11111011110110,
    14'b11111011111101,
    14'b11111100000011,
    14'b11111100000101,
    14'b11111100000101,
    14'b11111100000101,
    14'b11111100000101,
    14'b11111100001010,
    14'b11111100010010,
    14'b11111100011100,
    14'b11111100101100,
    14'b11111100111000,
    14'b11111101000011,
    14'b11111101001111,
    14'b11111101011111,
    14'b11111101101100,
    14'b11111101111000,
    14'b11111110001000,
    14'b11111110011100,
    14'b11111110101100,
    14'b11111110111011,
    14'b11111111001000,
    14'b11111111011100,
    14'b11111111101100,
    14'b11111111111000,
    14'b00000000001000,
    14'b00000000010010,
    14'b00000000010100,
    14'b00000000010111,
    14'b00000000010010,
    14'b00000000001101,
    14'b00000000000101,
    14'b11111111111011,
    14'b11111111101110,
    14'b11111111101110,
    14'b11111111110110,
    14'b00000000000000,
    14'b00000000010010,
    14'b00000000011111,
    14'b00000000100100,
    14'b00000000100100,
    14'b00000000011100,
    14'b00000000010100,
    14'b00000000001101,
    14'b00000000001000,
    14'b00000000010010,
    14'b00000000110001,
    14'b00000001010111,
    14'b00000010000101,
    14'b00000011000000,
    14'b00000100010100,
    14'b00000101001101,
    14'b00000101100110,
    14'b00000101100001,
    14'b00000100110001,
    14'b00000011101001,
    14'b00000010110001,
    14'b00000010000011,
    14'b00000001010010,
    14'b00000000001101,
    14'b11111111011100,
    14'b11111110111000,
    14'b11111110101001,
    14'b11111110110001,
    14'b11111111000101,
    14'b11111111011010,
    14'b11111111101100,
    14'b00000000000011,
    14'b00000000010111,
    14'b00000000101110,
    14'b00000000111101,
    14'b00000001001000,
    14'b00000001001111,
    14'b00000001001000,
    14'b00000000111101,
    14'b00000000101110,
    14'b00000000001101,
    14'b11111111111000,
    14'b11111111101001,
    14'b11111111011111,
    14'b11111111011100,
    14'b11111111100001,
    14'b11111111100100,
    14'b11111111100110,
    14'b11111111101001,
    14'b11111111101001,
    14'b11111111101100,
    14'b11111111101100,
    14'b11111111101110,
    14'b11111111101100,
    14'b11111111101100,
    14'b11111111101001,
    14'b11111111101110,
    14'b11111111110011,
    14'b11111111101110,
    14'b11111111101110,
    14'b11111111110011,
    14'b11111111110110,
    14'b00000000000000,
    14'b00000000001010,
    14'b00000000010100,
    14'b00000000100001,
    14'b00000000101100,
    14'b00000000110011,
    14'b00000000111000,
    14'b00000001000000,
    14'b00000001000011,
    14'b00000001001000,
    14'b00000001001010,
    14'b00000001001010,
    14'b00000001001010,
    14'b00000001001000,
    14'b00000001000000,
    14'b00000000110011,
    14'b00000000100100,
    14'b00000000011010,
    14'b00000000001101,
    14'b11111111101001,
    14'b11111111000101,
    14'b11111110110011,
    14'b11111110100110,
    14'b11111110011100,
    14'b11111110011010,
    14'b11111110000000,
    14'b11111101111011,
    14'b11111101100100,
    14'b11111101010010,
    14'b11111101001010,
    14'b11111101010100,
    14'b11111101101001,
    14'b11111110001010,
    14'b11111110011111,
    14'b11111110100110,
    14'b11111110100100,
    14'b11111110100001,
    14'b11111110100110,
    14'b11111110111000,
    14'b11111111001111,
    14'b11111111110110,
    14'b00000000001010,
    14'b00000000010111,
    14'b00000000100001,
    14'b00000000100110,
    14'b00000000100110,
    14'b00000000100110,
    14'b00000000100001,
    14'b00000000101001,
    14'b00000000011010,
    14'b00000000001000,
    14'b11111111100100,
    14'b11111110011010,
    14'b11111101010111,
    14'b11111100100100,
    14'b11111100001101,
    14'b11111101000011,
    14'b11111101100100,
    14'b11111110001010,
    14'b11111110101001,
    14'b11111111011010,
    14'b00000000000101,
    14'b00000000111101,
    14'b00000010000000,
    14'b00000011100110,
    14'b00000100101110,
    14'b00000101100110,
    14'b00000110001111,
    14'b00000110110011,
    14'b00000110111101,
    14'b00000110111101,
    14'b00000110101110,
    14'b00000110001101,
    14'b00000110000101,
    14'b00000101110011,
    14'b00000101100001,
    14'b00000101000101,
    14'b00000100101100,
    14'b00000100001111,
    14'b00000100000000,
    14'b00000011110011,
    14'b00000011101100,
    14'b00000011011111,
    14'b00000011001101,
    14'b00000010111011,
    14'b00000010110011,
    14'b00000010111011,
    14'b00000011001010,
    14'b00000011011100,
    14'b00000011101110,
    14'b00000011110011,
    14'b00000011101110,
    14'b00000011100001,
    14'b00000011001101,
    14'b00000010111011,
    14'b00000010101100,
    14'b00000010011100,
    14'b00000010001101,
    14'b00000001110011,
    14'b00000001011100,
    14'b00000001000000,
    14'b00000000100100,
    14'b11111111111101,
    14'b11111111101001,
    14'b11111111011010,
    14'b11111111010010,
    14'b11111111010100,
    14'b11111111011100,
    14'b11111111101100,
    14'b00000000001000,
    14'b00000000100100,
    14'b00000001000011,
    14'b00000001100001,
    14'b00000010001111,
    14'b00000010110011,
    14'b00000011010111,
    14'b00000100000000,
    14'b00000100111011,
    14'b00000101001101,
    14'b00000101010010,
    14'b00000101000000,
    14'b00000100101110,
    14'b00000100111011,
    14'b00000100110001,
    14'b00000101000101,
    14'b00000101001000,
    14'b00000101001101,
    14'b00000101011010,
    14'b00000101111000,
    14'b00000110101110,
    14'b00000111101110,
    14'b00001000001101,
    14'b00001000011111,
    14'b00001000011111,
    14'b00001000010010,
    14'b00001000000101,
    14'b00000111111101,
    14'b00000111111000,
    14'b00000111111011,
    14'b00000111110011,
    14'b00000111100110,
    14'b00000111001111,
    14'b00000110111000,
    14'b00000110001000,
    14'b00000101011111,
    14'b00000100110001,
    14'b00000100000101,
    14'b00000011010111,
    14'b00000010111000,
    14'b00000010100001,
    14'b00000010000101,
    14'b00000001100110,
    14'b00000001001101,
    14'b00000000111000,
    14'b00000000100110,
    14'b00000000010111,
    14'b00000000010100,
    14'b00000000011010,
    14'b00000000100001,
    14'b00000000100110,
    14'b00000000100001,
    14'b00000000011010,
    14'b00000000010100,
    14'b00000000010010,
    14'b00000000010010,
    14'b00000000010010,
    14'b00000000001111,
    14'b00000000001000,
    14'b11111111111011,
    14'b11111111110011,
    14'b11111111101100,
    14'b11111111101001,
    14'b11111111100100,
    14'b11111111100100,
    14'b11111111100100,
    14'b11111111100001,
    14'b11111111100100,
    14'b11111111101001,
    14'b11111111101110,
    14'b11111111110110,
    14'b11111111111101,
    14'b00000000000000,
    14'b00000000000011,
    14'b00000000000101,
    14'b00000000001000,
    14'b00000000001010,
    14'b00000000001010,
    14'b00000000001000,
    14'b00000000000101,
    14'b00000000000000,
    14'b11111111111101,
    14'b11111111111011,
    14'b11111111111000,
    14'b11111111110110,
    14'b11111111110011,
    14'b11111111110001,
    14'b11111111101110,
    14'b11111111101110,
    14'b11111111101110,
    14'b11111111110001,
    14'b11111111110011,
    14'b11111111110110,
    14'b11111111111000,
    14'b11111111111011,
    14'b11111111111101,
    14'b00000000000000,
    14'b00000000000000,
    14'b00000000000000,
    14'b00000000000011,
    14'b00000000000000,
    14'b00000000000000,
    14'b00000000000000,
    14'b11111111111101,
    14'b11111111111011,
    14'b11111111111011,
    14'b11111111111000,
    14'b11111111111000,
    14'b11111111110110,
    14'b11111111110110,
    14'b11111111110011,
    14'b11111111110110,
    14'b11111111110110,
    14'b11111111110110,
    14'b11111111111000,
    14'b11111111111000,
    14'b11111111111011,
    14'b11111111111011,
    14'b11111111111011,
    14'b11111111111101,
    14'b11111111111101,
    14'b11111111111101,
    14'b11111111111101,
    14'b11111111111101,
    14'b11111111111101,
    14'b11111111111101,
    14'b11111111111011,
    14'b11111111111011,
    14'b11111111111000,
    14'b11111111111000,
    14'b11111111110110,
    14'b11111111101100,
    14'b11111111011111,
    14'b11111111010111,
    14'b11111111011111,
    14'b11111111110011,
    14'b00000000010111,
    14'b00000000111011,
    14'b00000001010010,
    14'b00000001001010,
    14'b00000000101100,
    14'b00000000000101,
    14'b11111111100110,
    14'b11111111010100,
    14'b11111111011010,
    14'b11111111100100,
    14'b11111111101110,
    14'b11111111110001,
    14'b11111111101100,
    14'b11111111100110,
    14'b11111111100100,
    14'b11111111101001,
    14'b11111111110001,
    14'b11111111111101,
    14'b00000000000101,
    14'b00000000001010,
    14'b00000000001010,
    14'b00000000001000,
    14'b00000000000101,
    14'b00000000000011,
    14'b00000000000011,
    14'b00000000000101,
    14'b00000000001000,
    14'b00000000000011,
    14'b00000000000000,
    14'b11111111111011,
    14'b11111111110110,
    14'b11111111110001,
    14'b11111011111011,
    14'b11111000010111,
    14'b11110101100100,
    14'b11110111001000,
    14'b11111000100001,
    14'b11110111101100,
    14'b11110101111000,
    14'b11110101110011,
    14'b11110110010111,
    14'b11110111011111,
    14'b11111000100001,
    14'b11111000110011,
    14'b11111000101100,
    14'b11111000011010,
    14'b11111000010100,
    14'b11111000100110,
    14'b11111001011100,
    14'b11111011101100,
    14'b11111110000000,
    14'b00000001010100,
    14'b00000101001111,
    14'b00001001011010,
    14'b00001100001111,
    14'b00001101000011,
    14'b00001101010010,
    14'b00001101000000,
    14'b00001101010010,
    14'b00001101110110,
    14'b00001101111000,
    14'b00001101111000,
    14'b00001101011010,
    14'b00001011100100,
    14'b00001001011111,
    14'b00000111100100,
    14'b00000101101001,
    14'b00000011010010,
    14'b00000010000011,
    14'b00000001000101,
    14'b00000000000011,
    14'b11111110111000,
    14'b11111110000011,
    14'b11111101011100,
    14'b11111101010100,
    14'b11111101110011,
    14'b11111110100001,
    14'b11111111011010,
    14'b00000000100001,
    14'b00000001010010,
    14'b00000010000000,
    14'b00000010110001,
    14'b00000011100100,
    14'b00000100010010,
    14'b00000100101100,
    14'b00000011110011,
    14'b00000010110110,
    14'b00000001001000,
    14'b00000000010010,
    14'b11111111110011,
    14'b11111111101100,
    14'b11111111010111,
    14'b11111111000101,
    14'b11111110100100,
    14'b11111101111101,
    14'b11111101010100,
    14'b11111101001111,
    14'b11111101010100,
    14'b11111101100100,
    14'b11111110000011,
    14'b11111110010111,
    14'b11111110101110,
    14'b11111111001010,
    14'b11111111101100,
    14'b00000000001010,
    14'b00000000100110,
    14'b00000001000011,
    14'b00000001011111,
    14'b00000001101001,
    14'b00000001010111,
    14'b00000001000011,
    14'b00000000100100,
    14'b00000000010010,
    14'b00000000001101,
    14'b00000000001010,
    14'b00000000000101,
    14'b11111111110110,
    14'b11111111100110,
    14'b11111111010100,
    14'b11111111001000,
    14'b11111111000011,
    14'b11111111000011,
    14'b11111111001010,
    14'b11111111010010,
    14'b11111111011111,
    14'b11111111101001,
    14'b11111111110001,
    14'b11111111111101,
    14'b00000000001000,
    14'b00000000010010,
    14'b00000000011111,
    14'b00000000101100,
    14'b00000000101100,
    14'b00000000100100,
    14'b00000000010111,
    14'b00000000001101,
    14'b00000000001000,
    14'b00000000001010,
    14'b00000000001111,
    14'b00000000001010,
    14'b11111111110110,
    14'b11111111010100,
    14'b11111111001000,
    14'b11111111100001,
    14'b11111101010100,
    14'b11111001111000,
    14'b11110111100110,
    14'b11110101010111,
    14'b11111001001010,
    14'b11111011011100,
    14'b11111100100001,
    14'b11111011111011,
    14'b11111011101100,
    14'b11111100101110,
    14'b11111101111101,
    14'b11111111001000,
    14'b11111111110011,
    14'b11111111110001,
    14'b11111111000101,
    14'b11111110001101,
    14'b11111101001101,
    14'b11111100111000,
    14'b11111101001101,
    14'b11111101010111,
    14'b11111101000011,
    14'b11111101011010,
    14'b11111111010010,
    14'b00000010011111,
    14'b00000110111011,
    14'b00001001000000,
    14'b00001001011010,
    14'b00001000001000,
    14'b00000101001111,
    14'b00000011100001,
    14'b00000010110110,
    14'b00000011010100,
    14'b00000100011010,
    14'b00000101101100,
    14'b00000101111101,
    14'b00000101100100,
    14'b00000100110001,
    14'b00000011101100,
    14'b00000011001010,
    14'b00000010111000,
    14'b00000011000000,
    14'b00000011011100,
    14'b00000100001010,
    14'b00000100101001,
    14'b00000100111011,
    14'b00000101000101,
    14'b00000101001101,
    14'b00000101011100,
    14'b00000101111000,
    14'b00000110011100,
    14'b00000110111000,
    14'b00000111100110,
    14'b00001000001111,
    14'b00001000111000,
    14'b00001001011010,
    14'b00001001100110,
    14'b00001001100100,
    14'b00001001011100,
    14'b00001001001101,
    14'b00001000111011,
    14'b00001000100001,
    14'b00001000010010,
    14'b00001000000000,
    14'b00000111111000,
    14'b00000111111000,
    14'b00001000000000,
    14'b00001000000101,
    14'b00001000000000,
    14'b00000111110011,
    14'b00000111010111,
    14'b00000111001000,
    14'b00000111000000,
    14'b00000110111011,
    14'b00000110111011,
    14'b00000110110001,
    14'b00000101001111,
    14'b00000011001000,
    14'b00000000101001,
    14'b11111111111101,
    14'b00000000011111,
    14'b00000010000000,
    14'b00000011110110,
    14'b00000101110011,
    14'b00000111000011,
    14'b00001000001010,
    14'b00001001001010,
    14'b00001010010010,
    14'b00001011001000,
    14'b00001011100100,
    14'b00001011011111,
    14'b00001011011111,
    14'b00001011000101,
    14'b00001011011111,
    14'b00001100011111,
    14'b00001101101110,
    14'b00001110111000,
    14'b00001111000101,
    14'b00001110100110,
    14'b00001101111000,
    14'b00001100100110,
    14'b00001011101100,
    14'b00001010101100,
    14'b00001001110110,
    14'b00001000100110,
    14'b00000111100100,
    14'b00000110011111,
    14'b00000101011100,
    14'b00000011000000,
    14'b00000000011010,
    14'b11111100111000,
    14'b11111000100100,
    14'b11110010100110,
    14'b11101101110011,
    14'b11101100011100,
    14'b11110010000000,
    14'b11110111001010,
    14'b11111100101001,
    14'b00000010001111,
    14'b00000111001101,
    14'b00001011001010,
    14'b00001011111000,
    14'b00001011001101,
    14'b00001001011010,
    14'b00000111000101,
    14'b00000100001000,
    14'b00000010011111,
    14'b00000001110011,
    14'b00000001100110,
    14'b00000001010010,
    14'b00000000111011,
    14'b00000000100001,
    14'b00000000001010,
    14'b11111111110001,
    14'b11111111100100,
    14'b11111111111000,
    14'b00000000100001,
    14'b00000001011100,
    14'b00000010100100,
    14'b00000011011100,
    14'b00000100000101,
    14'b00000100101001,
    14'b00000101000011,
    14'b00000100110110,
    14'b00000100011100,
    14'b00000011111000,
    14'b00000011010010,
    14'b00000010011111,
    14'b00000010010010,
    14'b00000010010111,
    14'b00000010101110,
    14'b00000011000101,
    14'b00000011010111,
    14'b00000011001111,
    14'b00000011001000,
    14'b00000011000011,
    14'b00000011000101,
    14'b00000011000011,
    14'b00000010110011,
    14'b00000010001111,
    14'b00000001000000,
    14'b11111111110001,
    14'b11111110010111,
    14'b11111100110110,
    14'b11111011010100,
    14'b11111001010010,
    14'b11110111111000,
    14'b11110110101110,
    14'b11110101101100,
    14'b11110100100100,
    14'b11110100000000,
    14'b11110011101110,
    14'b11110011110001,
    14'b11110100010100,
    14'b11110101001101,
    14'b11110110010111,
    14'b11110111110011,
    14'b11111001111101,
    14'b11111011110011,
    14'b11111101100001,
    14'b11111110111011,
    14'b00000000001111,
    14'b00000000110110,
    14'b00000001001010,
    14'b00000001001111,
    14'b00000001001101,
    14'b00000001001000,
    14'b00000001000101,
    14'b00000001000000,
    14'b00000000111000,
    14'b00000000101001,
    14'b00000000011010,
    14'b00000000001101,
    14'b11111111111101,
    14'b11111111110001,
    14'b11111111011100,
    14'b11111111001101,
    14'b11111111000000,
    14'b11111110110110,
    14'b11111110100110,
    14'b11111110010111,
    14'b11111110001000,
    14'b11111101110001,
    14'b11111101000011,
    14'b11111100010010,
    14'b11111011100001,
    14'b11111010010100,
    14'b11111001011100,
    14'b11111000100110,
    14'b11110111110110,
    14'b11110110111101,
    14'b11110110101001,
    14'b11110110011010,
    14'b11110110001111,
    14'b11110110000101,
    14'b11110101111011,
    14'b11110110101110,
    14'b11110111001111,
    14'b11111000100100,
    14'b11111001101110,
    14'b11111010111011,
    14'b11111011101110,
    14'b11111100001010,
    14'b11111100001010,
    14'b11111011101110,
    14'b11111011000000,
    14'b11111010101110,
    14'b11111010101100,
    14'b11111010110011,
    14'b11111011000011,
    14'b11111011001010,
    14'b11111011010100,
    14'b11111011100001,
    14'b11111011101100,
    14'b11111011101110,
    14'b11111011110001,
    14'b11111011110110,
    14'b11111100000000,
    14'b11111100010010,
    14'b11111100101001,
    14'b11111101000101,
    14'b11111101110001,
    14'b11111110010111,
    14'b11111110111011,
    14'b11111111100001,
    14'b00000000000101,
    14'b00000000101110,
    14'b00000001010010,
    14'b00000010001111,
    14'b00000011000011,
    14'b00000011110001,
    14'b00000100011010,
    14'b00000101000000,
    14'b00000101101110,
    14'b00000110001000,
    14'b00000110011111,
    14'b00000110111011,
    14'b00000111010010,
    14'b00000111100110,
    14'b00000111111101,
    14'b00001000011100,
    14'b00001000111000,
    14'b00001001010100,
    14'b00001001010100,
    14'b00001001001000,
    14'b00001000101110,
    14'b00001000001111,
    14'b00001000001101,
    14'b00001000101110,
    14'b00001001101110,
    14'b00001011010100,
    14'b00001101011010,
    14'b00001101010010,
    14'b00001011011111,
    14'b00001001001000,
    14'b00000110110001,
    14'b00000011110011,
    14'b00000001111000,
    14'b00000000101001,
    14'b00000000010100,
    14'b00000000110110,
    14'b00000001011100,
    14'b00000001111011,
    14'b00000010010111,
    14'b00000010101110,
    14'b00000011001010,
    14'b00000011011100,
    14'b00000011110011,
    14'b00000100001111,
    14'b00000100111000,
    14'b00000101011010,
    14'b00000101110110,
    14'b00000110001010,
    14'b00000110011010,
    14'b00000110010100,
    14'b00000110000101,
    14'b00000101110011,
    14'b00000101011010,
    14'b00000101001101,
    14'b00000101001010,
    14'b00000101000000,
    14'b00000100111000,
    14'b00000101001101,
    14'b00000101010010,
    14'b00000101011010,
    14'b00000101100110,
    14'b00000101101001,
    14'b00000101100100,
    14'b00000101011111,
    14'b00000101011010,
    14'b00000101010111,
    14'b00000101011111,
    14'b00000101100100,
    14'b00000101101110,
    14'b00000101111011,
    14'b00000110001101,
    14'b00000110011111,
    14'b00000110110001,
    14'b00000111000011,
    14'b00000111001111,
    14'b00000111010111,
    14'b00000111011100,
    14'b00000111100110,
    14'b00000111110011,
    14'b00001000001000,
    14'b00001000010100,
    14'b00001000011111,
    14'b00001000100001,
    14'b00001000011111,
    14'b00001000001111,
    14'b00000111111101,
    14'b00000111100100,
    14'b00000111001010,
    14'b00000110101001,
    14'b00000110001111,
    14'b00000101111011,
    14'b00000101101001,
    14'b00000101010100,
    14'b00000101001000,
    14'b00000100111000,
    14'b00000100101110,
    14'b00000100100001,
    14'b00000100010111,
    14'b00000100001111,
    14'b00000100000101,
    14'b00000011111101,
    14'b00000011111011,
    14'b00000011111011,
    14'b00000011111000,
    14'b00000011111011,
    14'b00000011111011,
    14'b00000011111011,
    14'b00000011111011,
    14'b00000011111000,
    14'b00000011110001,
    14'b00000011100110,
    14'b00000011011010,
    14'b00000011001010,
    14'b00000010111000,
    14'b00000010100001,
    14'b00000010001111,
    14'b00000001111101,
    14'b00000001100100,
    14'b00000001000000,
    14'b00000000110011,
    14'b00000000010111,
    14'b11111111110011,
    14'b11111111001000,
    14'b11111110110001,
    14'b11111110011111,
    14'b11111110001000,
    14'b11111101111000,
    14'b11111101110001,
    14'b11111101101001,
    14'b11111101101001,
    14'b11111101011010,
    14'b11111101010010,
    14'b11111101001111,
    14'b11111101001111,
    14'b11111101001000,
    14'b11111100111000,
    14'b11111100011111,
    14'b11111100000101,
    14'b11111011100110,
    14'b11111010101100,
    14'b11111010000011,
    14'b11111001001111,
    14'b11111000101001,
    14'b11111000100110,
    14'b11111000111000,
    14'b11111001011111,
    14'b11111010010100,
    14'b11111100010010,
    14'b11111110101001,
    14'b00000001100100,
    14'b00000100101100,
    14'b00000110111011,
    14'b00000110110001,
    14'b00000110010111,
    14'b00000110101110,
    14'b00001000001111,
    14'b00001100000011,
    14'b00001110100100,
    14'b00001111101100,
    14'b00010000100100,
    14'b00010001000101,
    14'b00001111101001,
    14'b00001101010100,
    14'b00001011001111,
    14'b00001001101100,
    14'b00001000001111,
    14'b00000111000000,
    14'b00000110000011,
    14'b00000101000101,
    14'b00000011101001,
    14'b00000010101110,
    14'b00000001111101,
    14'b00000001010100,
    14'b00000000011100,
    14'b11111101000101,
    14'b11111100011010,
    14'b11111011111101,
    14'b11111100001000,
    14'b11111100111011,
    14'b11111110010111,
    14'b11111111110011,
    14'b00000001100100,
    14'b00000011000011,
    14'b00000100011111,
    14'b00000101101110,
    14'b00000110111101,
    14'b00000111000000,
    14'b00000110001000,
    14'b00000100101110,
    14'b00000010011100,
    14'b00000001010111,
    14'b00000000010111,
    14'b11111111001000,
    14'b11111110001101,
    14'b11111101111101,
    14'b11111101100001,
    14'b11111100011111,
    14'b11111101011111,
    14'b11111110100110,
    14'b11111110110110,
    14'b11111110110001,
    14'b11111111000011,
    14'b11111111011111,
    14'b00000000000000,
    14'b00000000010100,
    14'b00000000001111,
    14'b00000000011010,
    14'b00000000110001,
    14'b00000001000011,
    14'b00000001001000,
    14'b00000000101100,
    14'b11111111110110,
    14'b11111110101001,
    14'b11111101110011,
    14'b11111100111101,
    14'b11111100000101,
    14'b11111011011010,
    14'b11111010101100,
    14'b11111011000101,
    14'b11111011110001,
    14'b11111100000011,
    14'b11111011111011,
    14'b11111100001000,
    14'b11111100100001,
    14'b11111100110011,
    14'b11111100110110,
    14'b11111100110011,
    14'b11111100111000,
    14'b11111101000000,
    14'b11111101001000,
    14'b11111101001010,
    14'b11111101011010,
    14'b11111101111101,
    14'b00000001000000,
    14'b00000001111011,
    14'b00000010011100,
    14'b00000010110011,
    14'b00000010111011,
    14'b00000010110110
};

