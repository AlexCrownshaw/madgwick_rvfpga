`define ACC_WIDTH 11
`define ACC_INT_WIDTH 5
`define ACC_FRACT_WIDTH 6
`define GYRO_WIDTH 10
`define GYRO_INT_WIDTH 10
`define GYRO_FRACT_WIDTH 6
`define ACC_MAG_SQR_WIDTH 16
`define ACC_MAG_SQR_INT_WIDTH 12
`define ACC_MAG_SQR_FRACT_WIDTH 4
`define Q_HAT_DOT_MAG_SQR_WIDTH 16
`define Q_HAT_DOT_MAG_SQR_INT_WIDTH 12
`define Q_HAT_DOT_MAG_SQR_FRACT_WIDTH 4
`define Q_MAG_SQR_WIDTH 16
`define Q_MAG_SQR_INT_WIDTH 12
`define Q_MAG_SQR_FRACT_WIDTH 4
`define Q_WIDTH 16
`define Q_INT_WIDTH 2
`define Q_FRACT_WIDTH 14
`define Q_HALF_WIDTH 16
`define Q_HALF_INT_WIDTH 2
`define Q_HALF_FRACT_WIDTH 14
`define Q_TWO_WIDTH 17
`define Q_TWO_INT_WIDTH 3
`define Q_TWO_FRACT_WIDTH 14
`define Q_DOT_WIDTH 28
`define Q_DOT_INT_WIDTH 8
`define Q_DOT_FRACT_WIDTH 20
`define J_11_24_WIDTH 17
`define J_11_24_INT_WIDTH 3
`define J_11_24_FRACT_WIDTH 14
`define J_12_23_WIDTH 17
`define J_12_23_INT_WIDTH 3
`define J_12_23_FRACT_WIDTH 14
`define J_13_22_WIDTH 17
`define J_13_22_INT_WIDTH 3
`define J_13_22_FRACT_WIDTH 14
`define J_14_21_WIDTH 17
`define J_14_21_INT_WIDTH 3
`define J_14_21_FRACT_WIDTH 14
`define J_32_WIDTH 18
`define J_32_INT_WIDTH 4
`define J_32_FRACT_WIDTH 14
`define J_33_WIDTH 18
`define J_33_INT_WIDTH 4
`define J_33_FRACT_WIDTH 14
